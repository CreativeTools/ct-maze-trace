MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       ł���������������a������~g������~S�������j��������������~R������~b������~d�����Rich����                PE  L Gl�Q        � !
  v  �      �     �                       �                             �* K   % (                            p p  P�                            ` @            �                           .text   �t     v                   `.rdata  +�   �  �   z             @  @.data   |2   0                  @  �.reloc  �)   p  *   *             @  B                                                                                                                                                                                                                                                                                                                                                                                                V��> t�FP�7  ��V�7  ��^Ã�V�x7  ��^����U���E3��Y�   �A�A]� �����U��E�U�    �A�Q]� �������U����E�E���|�E�   ��C�H�U����   Vhp���    j3P��3����E�9u�~a�UJ�U�E�]��M��U  �M��[� �M�� t$ItIu0���K�@�D�����K�@�D�����K�@���U���F;u�|��E��M�jPQ�M��A  �E��+U����E�P�]��[6  �E���^��]�U���C�H���   ��$VWhp�jNj�ҋ}��������  �M��
��  �VUUU�����@S�]���M+UQPRW�}�E�����3�3��U܃��}�9M~L�E��� �Ut$HtHu2���S�@�T�����S�@�T�����S�@������AuGA;M|��}��C�؋H���   hp���    jiR�Ћ�C�Q���   �E�E+ǉE�hp���jjP��3Ƀ��E�9M~�U����E܉E�U��E����� �Ut(HtHu0���؋{�@�D�����؋{�@�D�����؋{�@�ǋ�������z�E�����E���E����E�A;M|�����E܋}�^�M�U�3��F�F�EP�E�GWQRPS�   �2����M�UQ�M�WR�F�E�PQS�����UR�F�\4  ��4[_��^��]ËE�~�F_�    ��^��]����������U���(SVW3����E������u�97��   �]��O�U�VUUU�����@��+�+�tHtHu�E���@��U���B��E��� �U��_����z
�O�E�   �u�U�ECSVR�UPR�n����E��g�E��������{�������A��   �}� �Ot�O�E�USVP�ERP�,��������   �E��   9w��   �]�G��M��4��E�H�v�$э��C�`�C�`������������������袗 �U�B�<� t'�M�����{�������Au��G�M����U���؋E�@�E�;G|���C�H�A�U�R�Ћ�C�Q�Jj j��E�hӑP�ыu����~|�	��$    ����C�B�P�M�Q�ҡ�C�H�Aj j��U�hБR�Ћ�C�Q�B<���M��Ћ�C�Q�RLj�j��M�QP�M��ҡ�C�H�A�U�R�Ѓ�Nu���C�Q�J�E�P�ыE���_^[��]� ��������������U���(��CS�]�CV�E�̑�Q���   hp���h�   P�ыs��3Ʌ�~��A;�|���C�E��B���   hp�jNj�у��E���@  �EW�}��U�Rj PV�'����U�3ۃ�3ɉ]��~"�U�R�}����@������AuCA;�|�]��C�؋Q���   hp���    jiP�ы�C��hp��E�B���   +���    jjQ���E؃�3҉E���~B�E��E�E�M����]�[�I������Au�E����E���E�����E�B;�|ʋ]�u�U�^�M�Qj3�R�F�F�E�S�]PS�   �����U�M�QjR�F�E�WPS������M�Q�F�:0  �U��4_�2^[��]ËM��H�M�p^�     �[��]��U��E� �M�������Au�ك����]� ������z	�   ]� 3�]� ���������  ��u��q  ��������������������������������U��E�� tHt	-�  3�]ùD��f  �����]ø   ]�����P�P��P(�P �P�P@�P8�P0�PX�PP�PH����������X�X�����������X�X �X(���������X0�X8�X@���XH���XP�XX��������U��M�U�A�
�E��B�I0���B�IH����A �
�A�A8�J���AP�J���X�A(�
�A�A@�J���AX�J���X�A�J�B �I0���B(�IH���X�A8�J �A �J���AP�J(���X �A@�J �A(�J���AX�J(���X(�A�J0�A0�J8���AH�J@���X0�A8�J8�A �J0���AP�J@���X8�A@�J8�A(�J0���AX�J@���X@�A�JH�BP�I0���BX�IH���XH�BP�I8�BH�I ���AP�JX���XP�A@�JP�BH�I(���AX�JX���XX]��̡�C�PH��p  j h�  Q�Ѓ�����̡�C�PH���   h�  Q�Ѓ��������U���C�HH���   SV�uWj h�  V�ҋء�C�HH���   h�  V�ҋM��3����s  �p���F�S(�<�    ��I �B��I �A�B��I8���B��IP���A(�J��A�A@�J����AX�J����B��I��B��I0���B��IH���Z����Z��Z��B��I �A�A8�J�����IP���B��I(�A�A@�J�����IX���B��I��B��I0����IH���Z����Z���A �J�A�B�I8���B�IP���A(�J�A�A@�J���AX�J���A�J��`N��B��I0���B��IH���Z����Z��Z��B��I �A�B��I8���AP�J����A(�J��A�B��I@���AX�J����B��I��B��I0���B��IH���Z����Z��Z�������u;�}j��T�+Ǎ�    �B���H�I �A�A8�J����B��IP���A(�J��A�A@�J����AX�J����B��I��B��I0���B��IH���Z����Z��Z�u���C���   �Bj j����_^[]� ��������U���C�H@�U�A,R�Ћ�C�Q��h�  �ȋB4h�  �и   ]� ������U���C�H�A��$�U�VR�Ћ�C�Q�Jj j��E�h �P�ы�C�B�P�M�Q�ҡ�C�H�Aj j��U�h�R�Ѓ�(�M�Q�M���i  � j P�U�Rh�0 jh'  �W  ��Ph�� �
q  ���M�����j  ��C�H�A�U�R�Ћ�C�Q�J�E�P�у���^��]�U���dS�]VW�M����]  ��C�HH���   S�҉E��C�PH�B$������P�MQ�U�R������U���   ���}��t(�MtQ�MpQ��`��R�U��   �M�R�|����   ��C�HH���   j S�҃���t&�Mt�UpQR��`��P�E�   �u�M�P�9����U��C�Q@�BS�Ѓ��   u<��C���   �Bh�  ���Ѕ�t �MpS��(  ��`���   �u�Mt�R  ��C���   �B4���Ћ؅�t=�Mt�Up�EQR��`���   �uS�M�P������C���   �B(���Ћ؅�u�_^[��]�p ���U���(  SV�M�W��h�����S  ��C���   �u�B4���Ћ�3�;�u3�_^[��]� �������]������jS�M�QjW�}W���k�  �E9]�uZ��C�BH���   WV�у��E�;�u=��C�BH���   jV�у��E�;�u��C�BH���   WV�у�_^[��]� S�u  ��C�B�P�M�Q�ҡ�C�H�ASj��U�h@�R�ЍM�Q�u  ��C�B�P�M�Q�ҡ�C�H@�Q,V�ҋ�C�Q��$h�  �ȋ��   h�  ��SP�E��e�  ���E�;�������M�Q�U�R��`�   ���E��E��E�   �������MPQ�M��]��]��]��]��]��]��]��]��]��]�������u��   ��P�����P�����`����5  V��P����  ��}��]�3��]��]ĉ]ԉ]̉]ȉ}�9]��  �]���U���4��]��C�HH���   h�  V�u��]��҃�����  �]����$    �u��C�HH��p  Sh�  V�ҋ���C�HH��p  }Sh�  V�ҋ�I�4ȋO�I�ЋO�&���C��|����f�I�C�E��f��� ���&�@�f�@�f���������������������������������������������R� ���8���E��]�9�|���th��E��&��C���f�C�f� �&�@�f�@�f���������������������������������������������߉ ���8��E��]�u��T����~��xjjjW���#  ��t	�F�E�����C�u܋QH�E����   �Eh�  FP�u��у�3�;��t����}��E�E��E����]�;�|jjjP�M���  ��t	�E�U���E�G�}�;}��������C�HH�u؋��   Sh�  V�҃�h�  ��h������CC  9]���  �E�;���  �}��E����$    ��h����5C  �M��]���E��|���S��4R��u�3ɉU���~*�E���������tA;�|���U��<��4I��u��M��ыE��؍�h����؍���B  ���C�QH��p  �]�j h�  W�Ћ�C�QH�؋��   h�  W�Ћ�C�QH��\�����   h�  W�Ћ�C�QH���   h�  W�E    ��H��$��~g�E��@�M�E�T����L��U���]�������C�HHt���   �Eh�  W��H��9E|����p  j h�  W�ҋ؋E����ء�C�HH��p  j h�  W�҃���h�������A  �]荍h����A  ݝx����K��S�M��h����E��U���A  �������z
�C9C��u�]�E��� ݅x������E��ʍ@�ǍǍ[���@���@������������� ���@���@�E��ˍ@������ ��ݝ8����@��ݝ@����@�E���݅8�����܅@������������������F����F0�����FH�����F ���F�F8�����FP�����F(�����F�F@�����FX����������Ƀ��M��X��E��X��S����u�3ۡ�C���   �BSj���Ћ�C���   �M�Bx�Ћ�C���   P�B|�����o  9]�t�M�Q�>!  ����P����]��]ĉ]ԉ]̉]��  9]�t�U�R�!  ���]��]��]��]��]�9]�t�E�P��   ��_��^[��]� �����U���VW�}���y
_3�^��]� S�]����  �F��;��ύ�N�U���u(��C�H��0  h��h@  �҃�[_3�^��]� ��;���  )^�F�Z  @����и   +�����ȋF�ڙ�ӉM�ȉE�ډU��������������]�;�u�;�u�;]�|�;M�r��]�Ù�E�9U��x���;��n����U�N�F�N��F��Ch����u�J�@���  ��hV  R�Ѓ���R�@hW  ��PQ��  �у��ȉ�������F�@�F��ʉN��~P+Ǎ@��P��+E�Í@��@�����R�P�� �N��+E��@����R�PQ�� ���  �@��+E����@��R�P�[�V  ��~�V�@���Q��RP謅 ���F�@���N�1  �F�D����@����E�F�ʙ�M�;���   	9E���   �E��������ً���������]�;������;������;]������	;M�������]�Ù�E�9U������;�������h����u$��C�H�E�@���  ��h{  R�Ѓ��$��C�Q�M�  �Ih|  ��QP�҃��ȉ���e����F�@����M�F�N�F;�})�N+Ǎ@�����R�P��@���R�h� ���} tA�N;�}��+��@�I��P��Nj Q較 ���[���R��Fj P衃 ���} tO�F;�}*�@��N��+ЉM�U��t������M��`�M�Mu�<��~��~��t��������`Ku�M��N[_�   ^��]� �����U���S�]V���y
^3�[��]� W�}���  �F��;��ˍ9�N�U���u(��C�H��0  h��h@  �҃�_^3�[��]� ��;��r  )~�F�8  @����и   +�������F�ʙ��߉}����ˋ�����ɉE����;�u��E�;�u�;�|�;�r��]�Ù9U�|�;�r��M�F�V��F�ы���Vh����u��C�Q���  hV  P�у����C�RhW  PQ��  �у���������V�}�N�ЉF��~B+��ɋ�+U��QӍЍQ��P�=� �F+]��    Q��RP�%� �����V  ��ɋ�+U�Q��Q��R�� ���3  ��~�V��    Q�R��R��� ���F����V�  �F�D����@����ȋF����M�;���   ;���   ������ɋ��;��6���;��.���;��&����}�;������E�;�����;������h����u#��C�Q���  ��    h{  P�у��"��C�Jh|  ��    RP��  �Ѓ����������N�]�ȉV�~�F;�}"�N�U+����P��P���Q�Ȁ ���} t?�F;�}�N��+����R��j R�� ���E�V��    Q��j P�� ���M��N_^�   [��]� ������������U��QSW��3�9tFV�w�]�9_~0��    9t	V�v  ���E���^�^�^�^@���E�;G|�W�P  ��^��_�_�_�__[��]���������U���S�]W��3�;����v���_�   [��]� V�w;�u(��C�H��0  h��h�  �҃�^_3�[��]� �G�D����@�ƙ���G�u��U�;�tG�w3ۉM�;�~59tV�  ��3ɃE���N�N�N�N�Gٙ��;�|�9E�rˋu��]�G��U�U��E�;�u	;U���   ;_~;U���   	;u���   �Ƌʋ�������������ɋ��;��4���;��,���;u��#����]�;������E�;��
���;�� ����h����u$��C�H���  �[���h�  R�Ѓ��$��C�Q��  �[��h�  �QP�҃��ȉ��������G�@���O�_�]3ɋG�[���RQP�} �E�O�3ۃ�3��]��E�;�|:;�v4�3�;�t�A   ��Y�Y�Y�Y�E���;�|��E�9E�r΋M^�O_�   [��]� �������Vh��jhPDj��  ������t���S  �,���^�3�^���������������U��S��V�s��y^3�[]�` jjjV������t�W�<v��{�   �u�_^�   []�` ����������U��M�U�A�
�E��A0�J���AH�J����A �
�A�A8�J���AP�J���X�A(�
�A�A@�J���AX�J���X]����U���C�HH���   SV�uWj h�  V�ҋء�C�HH���   h�  V�ҋM��3����s  �p���F�S(�<�    ��I �B��I �A�B��I8���B��IP���A(�J��A�A@�J����AX�J����B��I��B��I0���B��IH���Z����Z��Z��B��I �A�A8�J�����IP���B��I(�A�A@�J�����IX���B��I��B��I0����IH���Z����Z���A �J�A�B�I8���B�IP���A(�J�A�A@�J���AX�J���A�J��`N��B��I0���B��IH���Z����Z��Z��B��I �A�B��I8���AP�J����A(�J��A�B��I@���AX�J����B��I��B��I0���B��IH���Z����Z��Z�������u;�}j��T�+Ǎ�    �B���H�I �A�A8�J����B��IP���A(�J��A�A@�J����AX�J����B��I��B��I0���B��IH���Z����Z��Z�u���C���   �Bj j����_^[]� ��������U���C�H@�U�A,VR���X���C�QQ���$�B,h�  ���Ћ�C�Q�B0jh�  ���и   ^]� ���������U���C�H�A��$�U�VR�Ћ�C�Q�Jj j��E�h@�P�ы�C�B�P�M�Q�ҡ�C�H�Aj j��U�h8�R�Ѓ�(�M�Q�M��BR  � j P�U�Rh�F jh'  �@  ��Ph�� �jY  ���M����-S  ��C�H�A�U�R�Ћ�C�Q�J�E�P�у���^��]�U���|SV�uW�M�����  ��C�HH���   V�ҋء�C�PH�B$������P�MQ�U�R�6������   ���}��t'��`���E��P�   �MSQ�M������]��   ��C�BH�]���   j S�у���t%�U��`��RP�E�   �u�M�P�>����   ��C�Q@�BS�Ѓ��   uu��C���   �Bh$  ���Ѕ�tY��������ˋ�������~E���MQ�U�VR� �������̉�P�Q�P�Q�P�Q�P�@�Q�A�M�  ��Ou���C���   �B4���Ћ؅�t:���U��`���   �u�MQ�M�SR�p�����C���   �B(���Ћ؅�u�_^[��]�l ���������������U���  ��C���   �B4SV�u�M�W���Ћ�3�;���  �������]�����SS�M�QjW�}W��螐  ��C�E�BL�HxW�ы�C��h����B@�H,V���X���C�$���B���   h�  ����ݝ\�����C�P���   jh�  ���Љ�d���9]�u]��C�QH�u���   WV�Ѓ��E�;�u=��C�QH���   jV�Ѓ��E�;�u��C�QH���   WV�Ѓ�_^[��]� S�E�   �]��]��]��]��]��a]  ��C�Q�J�E�P�ы�C�B�PSj��M�h|�Q�ҍE�P�L]  ��C�Q�J�E�P�ыE��@���U�R�   �������M�u�PQ������j��\  ����h�  ����-  V�U�R�E�P����SS�E�   �]�]�]��]�]��n�  �����u�;�u<9]�t�M�Q�  ���]�]�]��]�]�9]�t�U�R�  ��3�_^[��]� �}�;���  �   W��l�����|�����l�����p����]���x�����t����	  W�M��u��]��]��]��]��]���  3��]�;�~��I ��p�����   @;�|�U����p������C�Q�J�E�P�]�ы�C�B�PSj��M�hh�Q�ҍE�P��[  ��C�Q�J�E�P���`��   �Ũ��U�;���  �E�Z   ����`��E��]��@�E�S�ЍM�Q�Mԍ�l���RP�E�P�2�������%  ��p������U����E�9�d���tZ���E�������A��   �E���������A�x   �E�����݅\�����������z^��������zY��+E�M�P�  �u�F݅\����]�����z6�E��E�;�|!jjjP�M��\  ��t�U�E���+M���u������ظgfff����������ɋ�+�u2�Eؙ����
P�RZ  ��h�����;�t��C�QPP�B�Ѓ���uv�ẼE�Z�]�F�E��]�;�������a��C�Q�J��T���P�ы�C�B�PSj���T���hH�Q�ҍ�T���P�Y  ��C�Q�J��T���P�у��~�������9}}%�u�;�|jjjV�M��X  ��t�E��+U���M��u�QW����t  ��C�BH���   Sh(  V�у�3�9]�~���    �U���ȉ\�A;M�|��C�HH���   Sh�  V�҃�3�;�~9�M����u��I�΋1�0�q�p�q�p�q�p�q�p�I�HB��;�|�9]�t�U�R��
  ���]��]��]��]��]�9�l���t��l���P��
  ���u܍M�Q��
  ��C���   �P��Sj���ҡ�C���   �M�Bx�Ћ�C���   P�B|�����<X  9]�t�M�Q�n
  ���]�]�]��]�]�9]�t�U�R�N
  ��_��^[��]� U���SVW�}3ۋ�;�)9t	V�"
  ��_��^�^�^�^^�   [��]� �N;�u(��C�H��0  h��h�  �҃�_^3�[��]� �F�D�����^@����E��U���t3�3Ʌ�~�Ù���� ;�|�;�r��}�F�M��;�u	9U���   ;�~9U���   ;���   �}����ɋ��;��z���;��r���;}��i����]�;��\����E�;��P���;��F����h����u#��C�Q���  ��    h�  P�у��"��C�Jh�  ��    RP��  �Ѓ����������N�}���V�^�N��    Pj Q��n �]�Ù��3�3Ʌ�|��t������ ;�|�;�r�_�^^�   [��]� ���������������U���VW�}���y
_3�^��]� S�]����  �F��;��ύ�N�U��u(��C�H��0  h��h@  �҃�[_3�^��]� ��;���  )^�F�b  @����и   +�����ȋF�ڙ�ӉM��ȉE��ډU����������ɋ���]�;�u�;�u�;]�|�;M�r��]�Ù�E�9U��u���;��k����U��N�F�N��F��Ch����u�J�@���  ���hV  R�Ѓ���R�@��hW  �PQ��  �у��ȉ��������F�@�F�щN��~P+Ǎ@���P��+E�Í@��P��@��P�m �N��ҋ�+E��R�@��RQ�gm ���  �@���P��+E��@��P�[�a  ��~�V����Q�R�@��R�!m ���F��@���V�7  �F�D����@����E��F�ʙ�M�;���   	9E���   �E���������ً�����ɋ���]�;������;������;]������	;M�������]�Ù�E�9U������;�������h����u'��C�H�E��@���  ���h{  R�Ѓ��'��C�Q�M���  �I��h|  �QP�҃��ȉ���Q����F�U��@���N�V�F;�}(�N+Ǎ@���P���P��@��P��k ���} tG�N;�}"��+��@���R�I�N��j R�(k ���V�[���P���j P�
k ���} tI�N��;�}�F�I�Ћ�+х�t�P�P���Ju�V��ʅ�~��t�P�P���Ku��؋E�F[_�   ^��]� ����U���S�]V���y
^3�[��]� W�}���  �F��;��ˍ9�N�U���u(��C�H��0  h��h@  �҃�_^3�[��]� ��;��j  )~�F�0  @����и   +�������F�ʙ��߉}����ˋ����ɉE����;�u��E�;�u�;�|�;�r��]�Ù9U�|�;�r��M�F�V��Fы���Vh����u��C�Q���  hV  P�у����C�RhW  PQ��  �у����� ����V�}�N���F��~@+�ɋ�+U��QӍ��Q��P�i �F+]��    Q��RP�i �����P  �ɋ�+U�Q��Q��R�zi ���/  ��~�V��    Q�R��R�Xi ���F����V�  �F�D����@����ȋF����M�;���   ;���   �����ɋ��;��@���;��8���;��0����}�;��#����E�;�����;������h����u#��C�Q���  ��    h{  P�у��"��C�Jh|  ��    RP��  �Ѓ����������N�]���V�~�F;�} �N�U+���P��P���Q�Dh ���} t=�F;�}�N��+���R��j R�g ���E�V��    Q��j P�g ���M��N_^�   [��]� ����������U��V���>  �Et	V�I  ����^]� ���������������Vh�jhPDj��  ������t���=  �N�d��,  ��^�3�^�������U��VW���w��y_3�^]� jjjV�.�����t�O�U�v����M�H�U�P�M�H�U�P�M_�H�   ^]� ���U��V��W�~��y_3�^]� jjjW�������t�F�M��_�   ^]� ������U��E��C� ]��U��V�u���t��C�QP��Ѓ��    ^]���������̡�C�H��@  hﾭ���Y����������U��E��t��C�QP��@  �Ѓ�]����������������U���C�H���  ]��������������U���C�H��  ]�������������̡�C�H��   ��U��E��t�x��u�   ]�3�]������U���s�   VW�xW�k ������u_^]Ã} tWj V�e ��_������F��C   ^]���U���C�E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�k ������u_^]�Wj V�d ��_������F��C   ^]�������������U���C�E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�j ������u_^]�Wj V�&d ��_������F��C   ^]�������������U���C�E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�j ������u_^]�Wj V�c ��_������F��C   ^]�������������U���C�E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�i ������u_^]�Wj V�&c ��_������F��C   ^]�������������U��M��t-�=�C t�y���A�uP��i ��]á�C�P�Q�Ѓ�]��������U��M��t-�=�C t�y���A�uP�i ��]á�C�P�Q�Ѓ�]��������U���C�H�U�R�Ѓ�]���������U���C�H�U�R�Ѓ�]���������U���C�E��t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   VW�xW�Vh ������u_^]�Wj V��a ��_������F��C   ^]���������U���C�E��tL�} t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   �U�IR�URP���  �Ѓ�]Ã�s�   VW�xW�g ������u_^]Ã} tWj V�3a ��_������F��C   ^]����������U��E��u�   ��C��t�U�IR�URP���   �Ѓ�]Ã�s�   VW�xW�'g ������u_^]�Wj V�` ��_������F��C   ^]����������U��E��u�   ��C��t,�} �U�IR�URPt���   �Ѓ�]Ë��  �Ѓ�]Ã�s�   VW�xW�f ������u_^]�Wj V� ` ��_������F��C   ^]�������U���C�H�U�R�Ѓ�]���������U���C�H�U�R�Ѓ�]���������U���C�H�U�R�Ѓ�]���������U���C�H�U�R�Ѓ�]���������U���C�Hp�]���C�Hp�h   �҃�������������U��V�u���t��C�QpP�B�Ѓ��    ^]���������U���C�Pp�EP�EPQ�J�у�]� U���C�Pp�EP�EPQ�J�у�]� U���C�Pp�EP�EPQ�J�у�]� U���C�Pp�EPQ�J�у�]� ����U��� �E�M���  �ȉESHV�u��W�}��A�Q����H։E��B��E���؉M�E��U���I �M��~�U�U�I)}�M��4�E��}���t�u+��\�P@�M���u�EH�E����   )}��u��	;]��u��s���u�]�;]}�M��>P�E�V�Ѕ�y�u�C�]�M��E��VP�҅��d����F��}��t�M�+���I ��P@�M��T�u�]��;]~��/���_^[��]� ������U���(W�}�����E�E�M���/  �ЉEH����B�J���SV�uƃ��ΉE��A��E����؉U��E܉M��
�U���$    ��~�M�M�J)}��U��G�M�E��M��t'�M�+����$    ��pf�\���M�f�f�4u�EH�E����   )}��u�;E��؉u�s���u�]�;]}�M��>P�E؋V�Ѕ�y�u�C�]��M��E�VP�҅��H����}�F���t!�M�+ȍI �Pf���Of�f�T�u�]��}�;E�~����	���^[_��]� ����������U���(W�}�����E�E�M���  �ЉEH����B�J���SV�uƃ��ΉE��A��E����؉U��E܉M��	�U���    ��~�M�M�J)}��U��9�M�E��M��t�M�+ȋ\�p���M��4u�EH�E����   )}��u�;E��؉u�s���u�]�;]}�M��>P�E؋V�Ѕ�y�u�C�]��M��E�VP�҅��W����}�F���t�M�+Ȑ��P��O��T�u�]��}�;E~��"���^[_��]� ��U��EP�u�E�UPR����]� 3҅��E�����UPRt	�+���]� �����]� ��������������U����ESV��W�]���t6�u��t/�}��t(�} t"�VP��Ѕ���   xO�E�   �}��}_^3�[��]� �}}���E������uu��VP�҅�tyO�}�G�}��E9E�~�_^3�[��]� ��~3�E���]��]�E����E�M���؋ESPO�҅�u����_��^[��]� �������U����ESV��W�]����  �u����   �}����   �} ��   �VP��Ѕ���   y�M_^�    3�[��]� �O�3��E�   �M��} ����   �EG�8_^3�[��]� �d$ �M�U���<�M������uuVQ���҅�ty�O��M��W�U��M9M�~�뤅�~1�E���]��]�E��E�M���؋ESPO�҅�u����_��^[��]� �M�9_^3�[��]� �U_^�����3�[��]� �������������U��V�u�F��F�����������������V ��������������D�Ez��^�P�P�]��������������N�X�N^�X]���������������U������P�M�P��P(�P �P�P@�P8�P0�PX�PP�XH���Q�P�Q�P�Q�P�Q�P�I�H�M��P�Q�P�Q�P �Q�P$�Q�P(�I�H,�M��P0�Q�P4�Q�P8�Q�P<�Q�P@�I�HD�M��PH�Q�PL�Q�PP�Q�PT�Q�PX�I�H\]� �����������U��y0 ts��U�����Au���A�Z����Au�B�Y�A�Z����Au�B�Y�A�����z��Y�A �Z����z�B�Y �A(�Z����zZ�B�Y(]� �E��Q�P�Q�P�Q �P�Q$�P�Q(�@�A,�Q�A��Q �A�A$�Q�Q(�A�A,�Q�A�A0   ]� U��V�u�������E���P�V�H�N�P�V�H�N�P�V��^]���������U��V�u���R����E� �^�@�^8�@���^X^]����������U���V�u�������E��_ �]��E��` �E��VX�������^@���^P�^8^��]�U���V�u���߿���E�_ �]��E�` �E��V�������^H���^(�^X^��]�U���V�u��蟿���E�W_ �]��E�|` �E��V�����V0���^ �^8^��]���U�������e�5���U��$�1a �m�����������E����������Az
���.���]��؋�]��������������U���h�E� V����u�������]����`�]��@�]�� �@�]��@�]���U����5���U��$�` �m�����������U��E����U����������Az�����]����]�������F���U��m����U��$�H` �m�����������U��E����U����������Az�����]����]�������F���U��m����U��$��_ �m�����������U��E����U����������Az�����]����]����������U��m����U��$�_ �m�����������U��E����U����������Az�����]����]�������F���U��m����U��$�J_ �m�����������U��E����U����������Az�����]����]�������F���U��m����U��$��^ �m��������^���E����������Az
������������E����E������������E����E������E�������������A�Eu�E���E��X�X��]����E���E��X�E��X��]�����������U�����V�u�V�VW�}��G����������fP �U����������Au>�����W��������z���_����^�^^��]����_����^�^^��]����_�������������z<��Az��������e�`�������u��������J����X �E������:��Az
������%�`�������u
���������X �E����������^ �^��_�^��^��]�U���PV�u�FP�M�Q�����FH�U����FP�]��FX�U����������7O �U����^������A��   �����U��E����E��E���������������Az�����)�`�������u
�����������5Y �E����������U�����z1�������������  �E��������E���X�X��]������������A�q  �E��������E���X�X��]����]����E�����������z<��Az��������e�`�������u��������J���$W �E������:��Az
������%�`�������u
����������V �E�������U���������Au����]�����}���\ �]��E��SY �]��E��xZ �E��M��E������������M�����������Az�����$�`�������u
���������W ���������]�����z�E���-���E��E���X�X��]ËE���E��E���X�X��]ËE���E���X�X��]������U���   V�u�������������Dz+�F��������Dz�F������Dz�u��螸����^��]�����U��{Y �]��E��@X ݝx����F�U��_Y �]��E��$X ݝp����F�U��CY �]��E��X �E����  �$�hc �E�u���E��E�P�ɍM�݅x���Q�ˍU�R�E���P�E��������������]������������]�݅p��������]������]������]��E����]������������]��������������]����]����U��U��]��[�����^��]��E��M���Q݅x����U���R�E��E���P�ˍM�Q�U��������]�݅p������E����������]������E������]��E��]������]��������]��������]������������]��  ���U��E�R�ɍE��E�P���M���Q�U�R�U������]��E���݅x��������]�݅p��������]������]������������]��E����������]������]������������]����  �E��E���P݅p����M���Q�E�U���R�ˍE�P�U�݅x��������E��������]������]��E����������]������������]��������]������������]����]��E����]����  �E�M���Q�E��U���R݅p����E���P�ʍM��E�Q�����������]������������]���݅x��������]������������]������������]��������]������]������]��E��   ���U��E�R�ɍE��E�P���M���Q�U�R�]�݅p������E��������]����]���݅x��������]������������]������]��������������]������E����������]��������]������������u�]�����U��U��]�������^��]Ð�_ �` !a �b �a .b U���xV�uW�   �}��E��P�M�Q�������H�U��P�M��H�U��P�@�M��M��U�Q�U�R�E�������P�M��H�U��P�M��H�UċP�EЉM�P�M�Q�U��~����E���E��H�UЋP�MԋH�U؋P�@�E�U��E������M����8���������u������`�������u
�������4R �}�u��EȍM��e�VQ��E��e��^�E��e��^��������H�N�P�V�H�N�P�V�@�F��������������Dz4�F��������Dz&�F��������Dz����������^�^�_^��]�_��^��]�������U���0V�uW�������}�������������Dz�G��������Dz�G��������D{�E����������Dz
_�؋�^��]��8��U��S �]��E��kR �]��E�WP������ �E������@���@�����Ȕ�������������E������]������]������������]��������������������������]��E����]����E������]��E��^�E��^ �E��^(�E������]��������������]����E�����_�]����E��^0�E��^8�E��^@���������������^H���^P�^X^��]����������������U��E�A    �]� �������������U��Q�@i�� %����E���E�y�ؔ�5Д��]�����U��Q�@i�� %����E���E�y�ؔ�5Д���%ؑ��]�������������U���V��~ ��   �Д�Ȕ������؋@i�� %����E��E�y�ؔ��@i�� ����%����U��E���E�y�ؔ�������U����������U�������t�����������D{�����������T ���u��D �E����F   �^^�M�����8���]��F�F    ���^�8���]������U���V��~ ��   �Д�Ȕ������؋@i�� %����E��E�y�ؔ��@i�� ����%����U��E���E�y�ؔ�������U����������U�������t�����������D{����������T ���u��C �E����F   �^^�M�����]��F�F    ��^��]��U��E�M�@�I�����A�H����� ���@�����H�E�������A�����X�i�X]�������U��E� ���@�@����������Au��������������Au����������������z��������������z����������������   ���������U�������z�E������������X�X��]���������������Dz�������+����������Dz���������Ȕ���������� ��5����������z
���ؑ�ɋE����E��X�X��]ËE�����������P�P���]������������U����E� �@�U��@�U�����������Au�E������������X�X��]�������������Dz����������U��$�HO �E����������E����E����������������������������5B H��wE�$�Lk �����ʋE��������X�X��]��������������ۋE��������X�X��]������k #k 'k +k /k U��M�A��A������������������������������Dz�E���P�P�]ËU�؋E�� �B�`�B�`������I���I����������I���I� �����@�@�E���������j�X�j�X]���̡�C�H���   ��U���C�H���   V�u�R�Ѓ��    ^]����������̡�C�H���   ��U���C�H���   V�u�R�Ѓ��    ^]����������̡�C�P���   Q��Y��������������U��� ��CSV��H�QPWV�u�����}�W�W3�����W(�E��W �_����_0����������_�_����������_���_ �_(;�~u��u���C�H�QLSV�ҋ����<t<uL�F(�E��f@P���]��F0�fH�]��F8�fP�]��i����F(�M��F@Q���]��FH�F0�]��F8�FP�]��C���C;]�|���_^[��]� ��U���C�P�EPQ���   �у�]� �U���C�P�EP�EP�EP�EP�EP�EPQ���   �у�]� �������������U���C�P�EP�EP�EP�EP�EP�EPQ���   �у�]� �������������U���C�P�EP�EP�EP�EPQ���   �у�]� �����U���C�P�EP�EP�EP�EPQ��  �у�]� �����U���C�P�EP�EP�EP�EPQ���  �у�]� �����U���C�P�EP�EPQ���   �у�]� �������������U��V�uW�����f  ��C�H���   VW�҃�_��^]� ��U���C�P�EPQ���   �у�]� �U���C�P�EPQ��  �у�]� ̡�C�P��0  Q�Ѓ�������������U���C�P�EP�EPQ��t  �у�]� �������������U���C�H�U���  j R�Ѓ�]���U���C�H���  V�u�R�Ѓ��    ^]�����������U���C�H���   ]��������������U���C�H���   V�u�R�Ѓ��    ^]�����������U��� ���C3��U�Q�U�Q�]�Q�M��M��P�E�PQ�E�P�EPPP�EP�EP�EP�EPQ��d  �у�8��]��������������U��U��tA���    t8��  �M;A}*V�1�0^t	�E�    �	��  �t	�E�    ]����U���C�H��P  ]��������������U���C�H��T  ]��������������U���C�H��X  ]�������������̋��     ��������V����t��C�QP��<  �Ѓ��    ^�����������U����t��C�Q�M���  Q�MQP�҃�]� ������U����t��C�Q�M���  Q�MQP�҃�]� ������U���C��S3�V��W�}��~D�^<�^8�^@�^H�FL   �^P�^T;���   �U�R���n  P�N诊  �M��7�  ���p  �F�E�P���x  ��N�P�V�H�N�P�V��C�H@�Q,W�ҋ���;�tG��C�P���   Sh6  ���ЉFP��C�Q���   Sh5  ����_�FT^[��]� �F   _^[��]� ���̋��@    � d   �V����t��C�QP��<  �Ѓ��    ^�����������U��V����t��C�QP��<  �Ѓ��    ��C�Q�E�MP�EQ��8  P��3҃����^��]� ���������U��E��u�D�MP�EPQ賤  ��]��������������̋�3ɉ�H�H�H�U��V��~ W�}u3h�j;hPDj��������t
W���N�  �3��F��u_^]� �~ t3�9_��^]� ��C�H<�W�҃�3Ʌ����_�F   ^��]� ��V���F   ��C�H<�Q��3Ʌ����^��������������̃y t�   ËA��uË�C�R<P��JP�у��������U����u��C�H�]� ��C�J<�URP�A�Ѓ�]� ���������������U��D��u��C�H�]Ë�C�J<�URP�A�Ѓ�]�U��D��$V��u��C�H�1���C�J<�URP�A�Ѓ�����C�Q�J�E�SP�ы�C�B�P�M�QV�ҡ�C�H�A�U�R�Ћ�C�Q�Jj j��E�hT�P�ы�C�B�@@�� j �M�Q�U�R�M��Ћ�C�Q�J���E�P���у���[t.��C�B�u�HV�ы�C�B�P�M�Q�҃���^��]á�C�P�E��RHjP�M��ҡ�C�P�E�M��RLj�j�PQ�M��ҡ�C�H�u�QV�ҡ�C�H�A�U�VR�Ћ�C�Q�J�E�P�у���^��]���������������U��D��$SV��u��C�H�1���C�J<�URP�A�Ѓ�����C�Q�J�E�P�ы�C�B�P�M�QV�ҡ�C�H�A�U�R�Ћ�C�Q�Jj j��E�hT�P�ы�C�B�@@�� j �M�Q�U�R�M��Ћ�C�Q�J���E�P���у���t/��C�B�u�HV�ы�C�B�P�M�Q�҃���^[��]á�C�P�E��RHjP�M��ҡ�C�P�E�M��RLj�j�PQ�M��ҡ�C�H�A�U�R�Ћ�C�Q�Jj j��E�hT�P�ы�C�B�@@��j �M�Q�U�R�M��Ћ�C�Q�J���E�P���у����3�����C�P�E��RHjP�M��ҡ�C�P�E�M��RLj�j�PQ�M��ҡ�C�H�u�QV�ҡ�C�H�A�U�VR�Ћ�C�Q�J�E�P�у���^[��]����������������U��D��$SV��u��C�H�1���C�J<�URP�A�Ѓ�����C�Q�J�E�P�ы�C�B�P�M�QV�ҡ�C�H�A�U�R�Ћ�C�Q�Jj j��E�hT�P�ы�C�B�@@�� j �M�Q�U�R�M��Ћ�C�Q�J���E�P���у���t/��C�B�u�HV�ы�C�B�P�M�Q�҃���^[��]á�C�P�E��RHjP�M��ҡ�C�P�E�M��RLj�j�PQ�M��ҡ�C�H�A�U�R�Ћ�C�Q�Jj j��E�hT�P�ы�C�B�@@��j �M�Q�U�R�M��Ћ�C�Q�J���E�P���у����3�����C�P�E��RHjP�M��ҡ�C�P�E�M��RLj�j�PQ�M��ҡ�C�H�A�U�R�Ћ�C�Q�Jj j��E�hT�P�ы�C�B�@@��j �M�Q�U�R�M��Ћ�C�Q�J���E�P���у����������C�P�E��RHjP�M��ҡ�C�P�E�M��RLj�j�PQ�M��ҡ�C�H�u�QV�ҡ�C�H�A�U�VR�Ћ�C�Q�J�E�P�у���^[��]��U��D��$SV��u��C�H�1���C�J<�URP�A�Ѓ�����C�Q�J�E�P�ы�C�B�P�M�QV�ҡ�C�H�A�U�R�Ћ�C�Q�Jj j��E�hT�P�ы�C�B�@@�� j �M�Q�U�R�M��Ћ�C�Q�J���E�P���у���t/��C�B�u�HV�ы�C�B�P�M�Q�҃���^[��]á�C�P�E��RHjP�M��ҡ�C�P�E�M��RLj�j�PQ�M��ҡ�C�H�A�U�R�Ћ�C�Q�Jj j��E�hT�P�ы�C�B�@@��j �M�Q�U�R�M��Ћ�C�Q�J���E�P���у����3�����C�P�E��RHjP�M��ҡ�C�P�E�M��RLj�j�PQ�M��ҡ�C�H�A�U�R�Ћ�C�Q�Jj j��E�hT�P�ы�C�B�@@��j �M�Q�U�R�M��Ћ�C�Q�J���E�P���у����������C�P�E��RHjP�M��ҡ�C�P�E�M��RLj�j�PQ�M��ҡ�C�H�A�U�R�Ћ�C�Q�Jj j��E�hT�P�ы�C�B�@@��j �M�Q�U�R�M��Ћ�C�Q�J���E�P���у����������C�P�E��RHjP�M��ҡ�C�P�E�M��RLj�j�PQ�M��ҡ�C�H�u�QV�ҡ�C�H�A�U�VR�Ћ�C�Q�J�E�P�у���^[��]����U���C�H<�A]����������������̡�C�H<�Q�����V��~ u>���t��C�Q<P�B�Ѓ��    W�~��t���z  W��������F    _^��������U���V�E�P���~�  ��P�������M���iz  ��^��]��̃=D uK�D��t��C�Q<P�B�Ѓ��D    �D��tV��� z  V�j������D    ^������������U���H��C�H�AS�U�V3�R�]��Ћ�C�Q�JSj��E�hX�P�ы�C�B<�P�M�Q�ҋ��C�H�A�U�R�Ѓ�;�u^3�[��]�V�M�]�蘪  �M�Q�U�R�M���  ���&  W�}�}���   ��C���   �U��ATR�Ћ�������   ��C�Q�J�E�P���ы�C�B���   ���M�Qj�U�R���Ћ�C�Q�J���E�P�ы�C�B�P�M�QV�ҡ�C�H�A�U�R�Ћ�C�Q�Bx��W�M����E���t�E� ��t��C�Q�J�E�P����у���t��C�B�P�M�Q����҃��}� u"�E�P�M�Q�M��ө  ��������E�_^[��]ËU��U�_�E�^[��]��U���DSV�u3ۉ]�;�u_��C�H�A�U�R�Ћ�C�Q�JSj��E�hX�P�ы�C�B<�P�M�Q�ҋ��C�H�A�U�R�Ѓ�;�u^3�[��]�V�M�]��Ѩ  �M�Q�U�R�M��!�  ���p  W�}��I �E����   ��C���   �U��ATR�Ћ�������   ��C�Q�J�E�P���ы�C�B���   ���M�Qj�U�R���Ћ�C�Q�J���E�P�ы�C�B�P�M�QV�ҡ�C�H�A�U�R�Ћ�C�Q�Bx��W�M����E��t�E ��t��C�Q�J�E�P����у���t��C�B�P�M�Q����҃��} tC�E�_^�E�[��]Ã�u1�E���t*��C���   P�BH�Ћ�C�Q���ȋBxW�Ѕ�t"�M�Q�U�R�M��§  ��������E�_^[��]ËM��M�_�E�^[��]�U��E��V3�;���   P�M��#�  �EP�M�Q�M�u��u�m�  ����   �u���E���tA��t<��uZ��C���   �M�PHQ�ҋ�C�Q���ȋBxV�Ѕ�u-�   ^��]Ë�C���   �E�JTP��VP�[�������uӍUR�E�P�M���  ��u�3�^��]����������V��~ u>���t��C�Q<P�B�Ѓ��    W�~��t���*u  W�t������F    _^�������̋�� h����������h����������̅�t��j�����̡�C�P��  ���C�P��(  ��U���C�P��   ��V�E�P�ҋuP���Zt  �M��t  ��^��]� ��������̡�C�P��$  ��U���C�H��  ]��������������U���C�H���  ]�������������̡�C�H��  ��U���C�H���  ]��������������U���C�H��x  ]��������������U���C�H��|  ]��������������U���EV���h�t	V���������^]� �������������̸   � ��������� ������������̸   � �������̸   � �������̸   � �������̸   � ��������� �������������3�� �����������3�� �����������3�� �����������3�� �����������3�� �����������3�� ����������̸   � �������̸   � �������̸   � ��������U���   V��诤  �����   �ESP�M���q  ��C�Q�J�E�P�ы�C�B�Pj j��M�hl�Q�҃��E�P�M��q  j j��M�Q�U�R��d���P��  ��P�M�Q�u  ��P�U�R�u  ���P�ϥ  ���M�����q  �M���q  ��d�����q  �M���q  ��C�H�A�U�R�Ѓ��M��q  ��[t	V�ߣ  ����^��]� ���U��EVP���a�  �����^]� �����Q誣  Y���������U��E�M�U�H4�M�P �U��M�@�� �@8�� �@<�� �@@�� �@D ��@H���@L@��@P0��@lP��@X�� �@\`� �@`���@d`��@T�� �@h���@pP� �@tp� �P0�H(�@,    ]��������������U���   h�   ��`���j P��$ �M�U�Ej Q�MRPQ��`���R�����E �Uh�   ��`���Q�E��ERPj�5  ��8��]��������������̋�`<����������̋�`0����������̋�`@����������̋�`����������̋�`����������̋�`����������̋�`����������̋�`,������������ �������������U���d�}W���*  ���Pt�U�S�U�]�]�S�҉E���  ��C�U�HH��   VRS�Ћ�C�Qd�J<�E��EP�эU�j/R���  �E�jP�  ��C�Qd�E�JpVSP�у�(3�j ��u��C�Bd�U�@�M�QR�����C�Qd�M�R�E�PQ��3���9u~b�3�;u���;�uO�E��RxVP�M�Q����� �U��@�]��@�]��������t��C�Hd�E���   j j�U�RP�у�F;u|�C���V���^[�   _��]� �������U����E�P�P�]� �������������  �������������3�� �����������U����   �ES��t
���[��]� ��C�PH�M�R,VW��$���P�ҋ���Pt�   �}��}W���E�����3��҅���   ���PxVW�M�Q����� �@�@���������A�|   �E���C�ˋUR�U��E����M����E������]��E����E��E������E������]��E������E��E������E������]�Hd�E�IP�ERP�у���t�E�u�t������؋�BtW��F��;��A����E�_^[��]� �����U�����CSVW�}��H@�Q8j W�ҋ]��Rx��SW�M�Q���ҋE�@��E�R|�Ƀ��ɋ�� �@0�E��������@H�E��������@ ���@�@8�����@P�����@(�����@�@@�����@X����S����������X�X�EP��_^�   [��]� ���������3�� �����������3�� ����������̸   �$ ��������� �������������� �������������� �������������3�� �����������3�� �����������U��UP�EQWRPV�<��������   ǆ�   p�ǆ�   ��ǆ�   �ǆ�   @� ǆ�   �� ǆ�   ��ǆ�    � ]������������U���C�P�B<��   V�u���Ѕ�t�Mj VQ��������u^��]�SWh   ������j R�C �]�E�}�M SP3��������(������E��� ��t�E�p� �� t�E�`� ��y�E�0� _��[t�E�P� �U�Eh   ������QRPj�b  ��^��]����������̋�`\����������̋�`l����������̋�`P����������̋�``����������̋�`p����������̋�`d����������̋�`X����������̋�`h�����������U���C�P8�EPQ�JD�у�]� ���̡�C�H8�Q<�����U���C�H8�A@V�u�R�Ѓ��    ^]�������������̡�C�H8�������U���C�H8�AV�u�R�Ѓ��    ^]��������������U���C�P8�EP�EP�EPQ�J�у�]� ������������U���C�P8�EP�EPQ�J�у�]� ��C�P8�BQ�Ѓ����������������U���C�P8�EPQ�J �у�]� ����U���C�P8�EP�EP�EP�EP�EPQ�J$�у�]� ����U���C�P8�EP�EP�EP�EP�EP�EPQ�J�у�]� U���C�P8�EP�EPQ�J(�у�]� U���C�P8�EP�EP�EPQ�J,�у�]� ������������U���C�P8�EP�EP�EPQ�J�у�]� ������������U���C�P8�EP�EP�EP�EP�EPQ�J�у�]� ����U���C�P8�EP�EPQ�J0�у�]� U���C�P8�EP�EP�EPQ�J4�у�]� ������������U���C�P8�EPQ�J8�у�]� ����U���C�H��x  ]��������������U���C�H��|  ]��������������U���C�H���  ]��������������U���C�H���  ]��������������U���C�H���  ]��������������U���C�H�A,]�����������������U���C�H�QV�uV�ҡ�C�H�Q8V�҃���^]�����̡�C�H�Q<�����U���C�H�I@]����������������̡�C�H�QD����̡�C�H�QH�����U���C�H�AL]�����������������U���C�H�IP]�����������������U���C�H��<  ]��������������U���C�H��,  ]��������������U���C�H�E���   �PPR�P@R�P0R�P R�PRP�EP�у�]������������̡�C�H���   ���C�H���  ��U���C�H�U�ER�UP�ER�UP���   Rh�.  �Ѓ�]����������������U���C�H�A]�����������������U���C�H��\  ]��������������U���C�H�AT]�����������������U���C�H�AX]�����������������U���C�H�A\]����������������̡�C�H�Q`����̡�C�H�Qd����̡�C�H�Qh�����U���C�H�Al]�����������������U���C�H�Ap]�����������������U���C�H�At]�����������������U���C�H��D  ]��������������U���C�H��  ]��������������U���C�H�Ix]�����������������U���C�H��@  ]��������������U��V�u���2b  ��C�H�U�A|VR�Ѓ���^]���������U���C�H���   ]��������������U���C�H��h  ]��������������U���C�H��d  ]��������������U���C�H���  ]�������������̡�C�H���   ��U���C�H��l  ]��������������U���C�H��   ]��������������U���C�H��  ]��������������U��V�u���>  ��C�H���   V�҃���^]���������̡�C�H��`  ��U���C�H��  ]��������������U���C�H�U���   ��R�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]�����U���C�H���  ]��������������U��U�E��C�H�E���   R���\$�E�$P�у�]�U���C�H���   ]��������������U���C�H���   ]��������������U���C�H���  ]��������������U���C�H���  ]��������������U���C�H���  ]��������������U���C�H���   ]��������������U���C�H���   ]��������������U���C�H���   ]��������������U���C�H���   ]��������������U���C�H���   ]��������������U���C�H���   ]��������������U�����C�P�E�P�E�P�E�PQ���   �у����#E���]����������������U�����C�P�E�P�E�P�E�PQ���   �у����#E���]����������������U�����C�P�E�P�E�P�E�PQ���   �у����#E���]����������������U���C�H��8  ]��������������U��V�u(V�u$�E�@��C�R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��V�u(V�u$�E�@��C�R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U���C�P0�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���   �у�(]�$ �U���C�P0�EP�EP�EP�EPQ���   �у�]� ����̡�C�P0���   Q�Ѓ�������������U���C�P0�EP�EPQ���   �у�]� �������������U���C�P0�EP�EP�EP�EPQ���   �у�]� ����̡�C�P0���   Q�Ѓ������������̡�C�H0���   ��U���C�H0���   V�u�R�Ѓ��    ^]�����������U���C�H��H  ]��������������U���C�H��T  ]�������������̡�C�H��p  ���C�H���  ��U���C�H���  ]��������������U���C�H���  ]��������������U���C�H���  ]��������������U���C�H���  ]��������������U���C�H���  ]��������������U���C�H�U�E��X  ��VR�UPR�E�P�ыu�    �F    ��C���   �Qj PV�ҡ�C���   ��U�R�Ѓ� ��^��]��������U���4VhLGOg�M��7  ��C�Q��X  3�VP�E�hicMCP�ы�C�u��u����   VP�A�U�R�Ћ�C���   �
�E�P�у� �M��r7  ��C���   �PT�M�Q�҃���u'�u����6  ��C���   ��U�R�Ѓ���^��]Ë�C���   �JT�E�P�ыu��P����6  ��C���   ��M�Q�҃���^��]���������������U���C�H��  ]��������������U���C�H��\  ]��������������U���C�H�U��t  ��V�uVR�E�P�у�����Z  �M���Y  ��^��]�����U���C�H�U���  ��VWR�E�P�ы�C�u���B�HV�ы�C�B�HVW�ы�C�B�P�M�Q�҃�_��^��]����������������U���C�H�U���  ��VWR�E�P�ы�C�u���B�HV�ы�C�B�HVW�ы�C�B�P�M�Q�҃�_��^��]����������������U���C�H���  ]��������������U���C�H���  ]��������������U���C�H���  ]��������������U���C�H���  ]��������������U���C�H���  ]��������������U���C�H�U�E��VWj R�UP�ERP��t  �U�R�Ћ�C�Q�u���BV�Ћ�C�Q�BVW�Ћ�C�Q�J�E�P�у�(_��^��]��U���C�H�U�E��VR�UP�ERP���  �U�R�Ћu�    �F    ��C���   j P�BV�Ћ�C���   �
�E�P�у�$��^��]���U���C�H��8  ]��������������U���  ��13ŉE��M�EPQ������h   R��b ����x	=�  |#���C�H��0  hp�hF  �҃��E� ��C�H��4  ������Rh���ЋM�3̓��D ��]�������U���C�H��  ��V�U�WR�Ћ�C�Q�u���BV�Ћ�C�Q�BVW�Ћ�C�Q�J�E�P�у�_��^��]����U���C�H��  ��V�U�WR�Ћ�C�Q�u���BV�Ћ�C�Q�BVW�Ћ�C�Q�J�E�P�у�_��^��]����U���C�H��p  ��4�҅���   h���M��%2  ��C�P�E�R4Ph���M��ҡ�C�P�E�R4Ph���M��ҡ�C�H��X  j �U�R�E�hicMCP�ы�C�E�    �E�    ���   j P�A�U�R�Ћ�C���   �
�E�P�ы�C���   ��M�Q�҃�$�M��1  ��]��������U���C�H��p  ��4V�҅�u��C�H�u�QV�҃���^��]�Wh!���M��,1  ��C�P�E�R4Ph!���M��ҡ�C�H��X  3�V�U�R�E�hicMCP�ы�C�u��u����   VP�A�U�R�Ћ�C���   �
�E�P�ы�C���   �PH�M�Q�ҋu����C�H�QV�ҡ�C�H�QVW�ҡ�C���   ��U�R�Ѓ�4�M��0  _��^��]������U���C�H��p  ��4V�҅�u��C�H�u�QV�҃���^��]�Wh����M��0  ��C�P�E�R4Ph����M��ҡ�C�H��X  3�V�U�R�E�hicMCP�ы�C�u��u����   VP�A�U�R�Ћ�C���   �
�E�P�ы�C���   �PH�M�Q�ҋu����C�H�QV�ҡ�C�H�QVW�ҡ�C���   ��U�R�Ѓ�4�M��/  _��^��]������U���C�H��p  ��4�҅�u��]�Vh#���M��$/  ��C�P�E�R4Ph#���M��ҡ�C�H��X  3�V�U�R�E�hicMCP�ы�C�u��u����   VP�A�U�R�Ћ�C���   �
�E�P�ы�C���   �P8�M�Q�ҋ��C���   ��U�R�Ѓ�(�M���.  ��^��]���������������U���C�H��p  ��4�҅�u��]�Vhs���M��D.  ��C�P�E�R4Phs���M��ҡ�C�H��X  3�V�U�R�E�hicMCP�ы�C�u��u����   VP�A�U�R�Ћ�C���   �
�E�P�ы�C���   �P8�M�Q�ҋ��C���   ��U�R�Ѓ�(�M���-  ��^��]���������������U���C�H���  ]��������������U���C�H��@  ]��������������U���C�H���  ]��������������U��V�u���t��C�QP��D  �Ѓ��    ^]������U���C�H��H  ]��������������U���C�H��L  ]��������������U���C�H��P  ]��������������U���C�H��T  ]��������������U���C�H��X  ]��������������U���C�H��\  ]�������������̡�C�H��d  ��U���C�H��h  ]��������������U���C�H��l  ]�������������̡�C�H���  ��U���C�H�U���  ��VR�E�P�ыu��P����+  �M���+  ��^��]�����U���C�H���  ]��������������U���C�H���  ]��������������U���C�H���  ]��������������U���C�H���  ]��������������U���C�H���  ]��������������U���C�H���  ]��������������U���C�H���  ]��������������U���C�H���  ]��������������U���C�H��$  ]��������������U���C�H��(  ]��������������U���C�H��,  ]�������������̡�C�H��0  ���C�H��<  ��U���C�H���  ]�������������̡�C�H���  ��U���C�H���  ]������������������������������U���C�H��  ]�������������̡�C�H��P  ���C���   ���   ��Q��Y��������U���C�H�A�U��� R�Ћ�C�Q�Jj j��E�h��P�ы�C�B�P�M�Q�ҡ�C�H�I�U�R�E�P�ы�C�B�P<�� �M��ҋ�C�Q�M�RLj�j�QP�M��ҡ�C�H�A�U�R�Ћ�C�Q�J�E�P�ы�C�B�P�M�Q�҃���]��������������U���C�E�PH�B���$Q�Ѓ�]� ���������������U���C�PH�EPQ���   �у�]� �U���C�PH�EPQ���  �у�]� �U���C�PH�EPQ���  �у�]� �U���C�PH�EP�EPQ��  �у�]� �������������U���C�PH�EP�EPQ��  �у�]� ������������̡�C�PH���  Q�Ѓ�������������U���C�PH�EPQ���  �у�]� ̡�C�PH���   j Q�Ѓ�����������U���C�PH�EPj Q���   �у�]� ��������������̡�C�PH���   jQ�Ѓ�����������U���C�PH�EPjQ���   �у�]� ��������������̡�C�PH���   jQ�Ѓ����������U���C�PH�EPjQ���   �у�]� ���������������U���C�PH�EP�EPQ���   �у�]� �������������U���C�PH�EP�EPQ���   �у�]� ������������̡�C�PH���   Q�Ѓ�������������U���C�PH�EP�EP�EP�EP�EPQ���  �у�]� �U��EVWP���@�  ������t�E��C�QH���   PVW�у���_^]� �����U��EVW���MPQ�L�  ������t�M��C�BH���   QVW�҃���_^]� ̡�C�PH���   Q�Ѓ������������̡�C�PH���   Q�Ѓ�������������U���C�PH�EPQ���   �у�]� �U���C�PH�EPQ���   �у�]� �U���C�PH�EP�EPQ��8  �у�]� �������������U���C�PH�EP�EPQ��   �у�]� ������������̡�C�PH���  Q�Ѓ������������̡�C�PH���  Q�Ѓ������������̡�C�PH���  Q�Ѓ������������̡�C�PH��  Q�Ѓ������������̡�C�PH��  Q�Ѓ�������������U���C�PH�EP�EPQ��  �у�]� �������������U���C�PH�EP�EP�EPQ��   �у�]� ���������U���C�PH�EP�EP�EP�EPQ��|  �у�]� �����U���C�PH�EPQ��  �у�]� ̡�C�PH��T  Q�Ѓ�������������U���C�PH�EP�EPQ��  �у�]� �������������U���C�PH�EPQ��8  �у�]� �U���C�PH�EPQ��<  �у�]� �U���C�PH�EPQ��@  �у�]� �U���C�PH�EP�EP�EPQ��D  �у�]� ��������̡�C�PH��L  Q��Y��������������U���C�PH�EPQ��H  �у�]� ̡�CV��H@�Q,WV�ҋ�C�Q��j �ȋ��   h�  �Ћ�C�QH�����   h�  V�Ѓ���
��t_3�^Ë�_^�̡�C�P@�B,Q�Ћ�C�Q��j �ȋ��   h�  �������U���C�E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U���C�E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U���C�PH�EP�EP�EPQ��   �у�]� ��������̡�C�HH��  ��U���C�HH��  ]��������������U���C�E�PH��$  ���$Q�Ѓ�]� �����������̡�C�PH��(  Q�Ѓ�������������U���C�PH�EP�EPQ��,  �у�]� �������������U���C�E�PH�EP�E���$PQ��0  �у�]� ���̡�C�PH���  Q�Ѓ������������̡�C�PH��4  Q�Ѓ������������̋��     �������̡�C�PH���|  jP�у���������U���C�UV��HH��x  R��3Ƀ������^��]� ��̡�C�PH���|  j P�у��������̡�C�PH��P  Q�Ѓ������������̡�C�PH��T  Q�Ѓ������������̡�C�PH��X  Q�Ѓ�������������U���C�PH��Q��\  �E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����̡�C�PH��`  Q�Ѓ�������������U���C�PH�EPQ��d  �у�]� �U���C�E�PH��h  ���$Q�Ѓ�]� ������������U���C�E�PH��t  ���$Q�Ѓ�]� ������������U���C�E�PH��l  ���$Q�Ѓ�]� ������������U���C�PH�EPQ��p  �у�]� �U���C�PH�EP�EP�EP�EPQ���  �у�]� �����U���C�PH�EP�EP�EP�EP�EP�EPQ���  �у�]� �������������U���C�E�HH�U �ER�UP�E���$R�UP���   R�Ѓ�]������������U��U�E��C�HH�E���   R�U���$P�ERP�у�]����������������U���E�M����  �M;�|�M;�~��]�����������U���C�PH�E���   Q�MPQ�҃�]� ������������̡�C�PH���   Q��Y�������������̡�C�PH���   Q�Ѓ������������̡�C�PH���   Q��Y��������������U���C�PH�EP�EPQ���   �у�]� �������������U���C�PH�EP�EP�EP�EP�EPQ���  �у�]� ̡�C�PH��t  Q��Y�������������̋�� ���@    ������C�Pl�A�JP��Y��������U���CV��Hl�V�AR�ЋE����u
�   ^]� ��C�Ql�MQ�MQ�
P�EP��3҃����F^��]� ������̋A��uË�C�QlP�B�Ѓ�������U���C�Pl�I�R�EP�EP�EP�EPQ�ҋE�M��;�u�E]� 9Mt���]� ������������U��U�E��C�HH�ER�U���$P���  R�Ѓ�]����U���C�HH���  ]��������������U���C�HH���  ]��������������U��U0�E(��C�HH�E$R�U ���$P�ER�UP�ER�UP�ER�UP���  R�Ѓ�,]������������U���C�HH���  ]��������������U���C�E�PH�EP���$Q���  �у�]� ��������U���SV��豈  �؉]����   �} ��   ��C�HH��p  j h�  V�҃��E��u
^��[��]� �MW3��}����  ����   �]��I �E�P�M�Q�MW��  ��t_�u�;u�W�I ������u�E����ҋL�;L�t-��C�Bl�S�@����QR�ЋD������t	�M�P�e�  F;u�~��}��MG�}��0�  ;��x����]�_^��[��]� ^3�[��]� U�����CSV�ًHH��p  j h�  S�]��ҋ�����u
^3�[��]� �E��u��C�HH���  �'��u��C�HH���  ���uš�C�HH���  S�ҋȃ��E��t�W��  ��C�HH���   h�  S3��҃����  ���_�u����    ��C�Hl�U�B�IWP�ы�������   ��C�F�J\�UP�A,R�Ѓ���t�K�Q�M�%�  ��C�F�J\�UP�A,R�Ѓ���t�K�Q�M���  �E��;Pt&�F��C�Q\�J,P�EP�у���t	�MS�̆  ��C�v�B\�M�P,VQ�҃���t�M�CP裆  ��C�QH�E����   �E�h�  PG���у�;�����_^�   [��]� ��������U���C�HH���   ]�������������̡�C�PH���   Q��Y��������������U���C�HH���  ]��������������U���C��P���   V�uW�}���$V�����E������At���E������z����؋�C�Q�B,���$V����_^]����������������U���0���C�U�V�u�U��]�W�P�}���   �E�PV�M�Q����� �@�@�E�����E��Au�����������z���������������z�����������Au������������z)���١�C�]��ɋ��]��]��P�RH�E�PV��_^��]���������Au������������������U���C�HH�]��U���C�H@�AV�u�R�Ѓ��    ^]�������������̡�C�HH�h�  �҃�������������U���C�H@�AV�u�R�Ѓ��    ^]��������������U���C�HH�Vh  �ҋ�������   �EPh�  �~  ����t]��C�QHj P���   V�ЋMQh(  �f~  ����t3��C�JH���   j PV�ҡ�C���   �B��j j���Ћ�^]á�C�H@�QV�҃�3�^]�������U���C�H@�AV�u�R�Ѓ��    ^]��������������U���C�HH�Vh�  �ҋ�����u^]á�C�HH�U�E��  RPV�у���u��C�B@�HV�у�3���^]�������U���C�H@�AV�u�R�Ѓ��    ^]��������������U���C�HH�I]�����������������U���C�H@�AV�u�R�Ѓ��    ^]��������������U���C�PH�EPQ���  �у�]� �U���C�PH�EPQ���  �у�]� ̡�C�PH���  Q�Ѓ�������������U���C�HH���  ]��������������U���C�E�HH�U0�E,R�U(P�E$R�U P�ER�U���\$�E�$P��P  R�Ѓ�,]������������̡�C�PH���  Q�Ѓ�������������U���C�PH�EP�EPQ���  �у�]� ������������̡�C�PH��  Q�Ѓ�������������U���C�PH�EP�EP�EPQ���  �у�]� ��������̡�C�PH���  Q�Ѓ������������̡�C�PH���  Q�Ѓ�������������U���C�PH�EPQ��  �у�]� �U���C�PH�EPQ��  �у�]� ̋������������������������������̡�C�HH���  ��U���C�HH���  ]��������������U���C�PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ���������U���C�PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ��������̡�C�PH��,  Q�Ѓ�������������U���C�PH�EPQ��X  �у�]� ̡�C�PH��\  Q�Ѓ�������������U���C�HH��0  ]��������������U���C��W���HH���   j h�  W�҃��} u�   _��]� Vh�  �y  ��������   ��C�HH���   j VW�҃��M��C  ��C�P�E�R0Ph�  �M����E��C�P�B,���$h�  �M��Ћ�C�Q@�J(j �E�PV�у��M��L  ^�   _��]� ^3�_��]� �����U��S�]�; VW��u7��C�U�HH���   RW�Ѓ���u��C�QH���   jW�Ѓ���t�   �����   ��C�QH���   W�Ѓ��} u(��C�E�QH�M���  P�ESQ�MPQW�҃��B�u��t;��C�U�HH�ER�USP���  VRW�Ћ�C���   �B(�����Ћ���uŃ; u��C�QH���   W�Ѓ���t3���   �W��u1��C�QH���   �Ћ�C�E�QH���   PW�у�_^[]� ��C�BH���   �у��} u0��C�M�BH�U���  Q�Mj R�UQRW�Ѓ�_^��[]� ��C�QH�h  �Ћ؃���u_^[]� ��C���   �u�Bx���Ћ�C���   P�B|���Ѕ�tU��C�E�QH�MP�Ej Q���  VPW�у���t��C���   �ȋBHS�Ћ�C���   �B(���Ћ���u�_^��[]� ��������������U��EV���u��C�HH���  �'��u��C�HH���  ���u��C�HH���  V�҃���u3�^]� P�EP���N���^]� ���������U���D��C�HH���   S�]VWh�  S�ҋ��C�HH���   3�Wh�  S�u܉}��҃��E�}�}��}�;��>
  ��C���   �B���Ћ�C=�  �  �QH���   Wh:  S�Ћ�C�QH�E����   h�  S�Ћ�C�QHW�����   h�  S�uԉ}��Ћ�C�QH�E苂  S�Ћ�C�QH�EЋ��  S�Ѓ�(�E��E�̕��~~�M���M�I �MЅ�tMj�W豋  ���t@�@�Ẽ|� �4�~����%�������;�u/���0�  ;E�~�E؋���  E���E�;Pu�E���E��E�G;}�|��}� ��   �u�j S���t  ����  ���Xw  ��ti���q  �}�;�u^��C�H���  �4�hЕ��h�  V�҃��E���b  �M��E��	w  ��t�}� t��tVP�E�P�p�  ����}܋�C�Q���  �4�hЕ��h�  V�Ѓ��E����  �M�3�;�t;�tVQP� �  ���E�;�~-��C�QhЕ��h�  P���   �Ѓ��E�;���  ��C�E��QH��  j�PS�у�����  �u�;�tjS����r  ���{  ���Fv  �E���}��C�BH���   Wh�  S�у�3��E�}�9}��]  �}���}����$    �MЅ��J  �U�j�R蚉  ����6  �M̍@�|� ���]�~����%�������9E���  ���ݒ  �E�3�3ɉE܉M�9C��   ��$    �����������ti�]������������M�ҋ9�<��}�҉T��y�]��|��]��z�|��y�]��|��]��z�|��I�}��]��L��M��}ȃ��T����M�A�M�;K�v����E؅��0  �+U�j��PR�M��W����M�v���E�3�+��U��E��ʋE�;E���   �}� �U����E�t4�U�M��@���P�Q�P�Q�P�Q�P�Q�@�A�M��Eȍ@�E��Ћ��P�Q�P�Q�P�Q�P�Q�@�A;]�}_�UȋE�9�uT�ȋL�����������w0�$�$� �U���4���M���t���U���t��	�M���t��M���;]�|��E܃�F�M�;]������U�;U��  �U�R��w���E�P��w���M�Q�w����_^3�[��]Ë�M�3�;G�Å���   �E�v�ЋW��R�ы��Q�P�Q�P�Q�P�Q�P�I�H�O��I�M�ы�P�Q�P�Q�P �Q�P$�Q�P(�I�H,��@�E�ЋU�Lv�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��t8�G�U�@�ʋU�Lv	�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��w��U��@�ʋU�F�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��w��U�F�@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�7F��t=�G�U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�wF���O�E�@���E��}�;E�������U�R�u���E�P�u�����  ���   �B����=  ��  ��C�QH���   j h(  S�Ћ�C�QH�����   h(  S�ЋЃ�3��U؅�~"��ǅ�t�|� t�4N��tN�@;�|�u��u܋�C�Q���  �4v�hЕ��hK  V�Ѓ��E�����   �M��t��tVQP�8�  ���u؋�C�Q���  �hЕ��hP  V�Ѓ��E���tP��t��tVWP���  ���M����+�C�RH��PQ�E���   S�Ѓ���u�M�Q�bt���U�R�Yt����_^3�[��]á�C�HH���   j h�  S�҉E���C�HH���   j h(  S��3�3���3��E��}ĉ]�9]��:  �U��څ��  �E�    ����   �U�<��v��   ����U��:��\:�Y�\:�Y�\:׉Y�Z�Y�R�Q�U��\�EԉY�\�T�Y�Z�Y �Z�Y$�Z�Y(�R�]��Q,�U�@����0��;�|��}ă|� �t   �U��M�ύI�ʋU�v���A�B�A�B�A�B�A�B�I�J�E���ЋE�Tv�Ћ��A�B�A�B�A�B�A�B�I�J�U���<ډ}�C�]�;]�������M�3�3�;�~�U���$    �t���   @;�|��U�R�r�����E�P�r����_^�   [��]�{� �� �� �� ������������U��E� �M+]� ���������������U��V��V�����C�Hl�AR�Ѓ��Et	V�Tu������^]� ���������̡�C�P�BVj j����Ћ�^���������U���C�P�E�RVj P���ҋ�^]� U���C�P�E�RVPj����ҋ�^]� ��C�P�B�����U���C�P���   Vj ��Mj V�Ћ�^]� �����������U���C�P�EPQ�J�у�]� ����U���C�P�EPQ�J�у����@]� ���������������U���C�P�E�RtP�ҋ�C���   P�BX�Ѓ�]� ���U���C�P�E�Rlh#  P�EP��]� ���������������U���C�P�E�RlhF  P�EP��]� ���������������U���C�P�E�RtP�ҋ�C���   �M�R`QP�҃�]� ���������������U���C�P���   ]��������������U���C�P�E���   P�҅�u]� ��C���   P�B�Ѓ�]� �������̡�C�HL���   ��U���C�H@�AV�u�R�Ѓ��    ^]�������������̡�C�HL�������U���C�H@�AV�u�R�Ѓ��    ^]�������������̡�C�PL���   Q�Ѓ�������������U���C�PL�EP�EPQ���   �у�]� �������������U���CV��HL���   V�҃���u��C�U�HL���   j RV�Ѓ�^]� ��C���   �ȋBP�Ћ�C���   �MP�BH��^]� �����̡�C�PL��(  Q�Ѓ�������������U���C�PL�EP�EPQ��,  �у�]� ������������̡�C�HL�Q�����U���C�H@�AV�u�R�Ѓ��    ^]��������������U���C�PL�E�R��VPQ�M�Q�ҋu��P���%����M��=�����^��]� ����U���C�PL�EPQ���   �у�]� �U���C�PL�EP�EPQ�J�у�]� ��C�PL�BQ�Ѓ���������������̡�C�PL�BQ�Ѓ���������������̡�C�PL�BQ�Ѓ����������������U���C�PL�EP�EP�EPQ�J �у�]� ������������U���C�PL�EPQ��4  �у�]� �U���C�PL�EP�EP�EPQ�J$�у�]� ������������U���C�PL�EP�EP�EP�EPQ�J(�у�]� �������̡�C�PL�B,Q�Ѓ���������������̡�C�PL�B0Q�Ѓ����������������U���C�PL�EP�EPQ��  �у�]� ������������̡�C�PL���   Q�Ѓ�������������U���C�PL�E��  ��VPQ�M�Q�ҋu��P�������M�������^��]� ̡�C�PL�B4Q�Ѓ���������������̡�C�PL�B8j Q�Ѓ��������������U���C�PL���   ]��������������U���C�PL���   ]��������������U���C�PL���   ]��������������U���C�PL���   ]��������������U���C�PL���   ]��������������U���C�PL���   ]��������������U���C�PL���   ]��������������U���C�PL���   ]��������������U���C�PL���   ]��������������U���C�PL�EPQ�J<�у�]� ���̡�C�PL�BQ��Y�U���C�PL�EP�EPQ�J@�у�]� U���C�PL�Ej PQ�JD�у�]� ��U���C�PL�Ej PQ�JH�у�]� ��U���C�PL�EjPQ�JD�у�]� ��U���C�PL�EjPQ�JH�у�]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}���G  W�M�Q�U�R���č  ���M����W:  ��t��C���   ��U�R�Ѓ�_^3�[��]Ë�C���   �J8�E�P�ы�C�����   ��M�Q�҃�_��^[��]��������������U���$3�V�E��E�E��P�M��E�   �E�   �E��  �>G  j�M�Q�U�R���-�  �M��9  ��C���   ��U�R�Ѓ�^��]�����������U���$��C�UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}��F  j�E�P�M�Q��詌  �M��!9  ��C���   ��M�Q�҃�_^��]� ��U���$��C�UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}��:F  j�E�P�M�Q���)�  �M��8  ��C���   ��M�Q�҃�_^��]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}���E  W�M�Q�U�R��褋  ���M����78  ��t+�u���	  ��C���   ��U�R�Ѓ�_��^[��]� ��C���   �JL�E�P�ыu��P���u  ��C���   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}��E  W�M�Q�U�R����  ���M����w7  ��t+�u���I  ��C���   ��U�R�Ѓ�_��^[��]� ��C���   �JL�E�P�ыu��P���  ��C���   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}��TD  W�M�Q�U�R���$�  ���M����6  _^��[t��C���   ��U�R�������]Ë�C���   �J<�E�P���]���C���   ��M�Q���E�����]���������������U���$SVW3��E��P�M��}܉}��E��  �}��}��C  W�M�Q�U�R���t�  ���M����6  ��t��C���   ��U�R�Ѓ�_^3�[��]Ë�C���   �J8�E�P�ы�C�����   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}���B  W�M�Q�U�R���Ĉ  ���M����W5  ��t-��u��C����   ���^�U�R�Ѓ�_��^[��]� ��C���   �JP�E�P�ы�u�H��P�@�N��C�V���   �
�F�E�P�у�_��^[��]� �����̡�C�PL���   Q��Y��������������U���C�PL�E���   ��jPQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U���C�PL�E���   ��j PQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U���$SVW3��E��P�M��}܉}��E��  �}��}��dA  W�M�Q�U�R���4�  ���M�����3  ��t-��u��C����   ���^�U�R�Ѓ�_��^[��]� ��C���   �JP�E�P�ы�u�H��P�@�N��C�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��@  W�M�Q�U�R���d�  ���M�����2  ��t-��u��C����   ���^�U�R�Ѓ�_��^[��]� ��C���   �JP�E�P�ы�u�H��P�@�N��C�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}���?  W�M�Q�U�R��蔅  ���M����'2  ��t-��u��C����   ���^�U�R�Ѓ�_��^[��]� ��C���   �JP�E�P�ы�u�H��P�@�N��C�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}���>  W�M�Q�U�R���Ą  ���M����W1  ��t��C���   ��U�R�Ѓ�_^3�[��]Ë�C���   �J8�E�P�ы�C�����   ��M�Q�҃�_��^[��]��������������U����E3�V�]�E��E��E��P�M�E�   �E��  �?>  j�M�Q�UR���.�  �M�0  ��C���   ��U�R�Ѓ�^��]� ���������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E���=  j�U�R�E�P��较  �M��60  ��C���   �
�E�P�у�^��]� ��������U���$��C�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��J=  j�E�P�M�Q���9�  �M��/  ��C���   ��M�Q�҃�_^��]� ��U���$��C�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}���<  j�E�P�M�Q��蹂  �M��1/  ��C���   ��M�Q�҃�_^��]� ��U���$��C�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��J<  j�E�P�M�Q���9�  �M��.  ��C���   ��M�Q�҃�_^��]� ��U���$��C�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}���;  j�E�P�M�Q��蹁  �M��1.  ��C���   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��_;  j�U�R�E�P���N�  �M���-  ��C���   �
�E�P�у�^��]� ��������U���$SVW3��E��P�M��}܉}��E��  �}��}���:  W�M�Q�U�R���Ā  ���M����W-  ��t-��u��C����   ���^�U�R�Ѓ�_��^[��]� ��C���   �JP�E�P�ы�u�H��P�@�N��C�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��$:  W�M�Q�U�R����  ���M����,  ��t��C���   ��U�R�Ѓ�_^3�[��]Ë�C���   �J8�E�P�ы�C�����   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}��t9  W�M�Q�U�R���D  ���M�����+  ��t��C���   ��U�R�Ѓ�_^3�[��]Ë�C���   �J8�E�P�ы�C�����   ��M�Q�҃�_��^[��]��������������������t��t��t3�ø   ����U���$��C�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��8  j�E�P�M�Q���y~  �M���*  ��C���   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��8  j�U�R�E�P���~  �M��*  ��C���   �
�E�P�у�^��]� ��������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��7  j�U�R�E�P���}  �M��*  ��C���   �
�E�P�у�^��]� ��������U���C�H���   ]��������������U���C�H���   ]�������������̡�C�H���   ���C�H���   ��U���C�H���   V�u�R�Ѓ��    ^]�����������U���C�H���   ]��������������U���C�HL�QV�ҋ���u^]á�C�H�U�ER�UP���  RV�Ѓ���u��C�Q@�BV�Ѓ�3���^]����������U���C�H�U�E���  R�U�� P�ERP�у�]������U���C�H���   ]��������������U���C�H�U �ER�UP�ER�UP�ER�UP���   R�Ѓ�]������������̡�C�PL�BLQ�Ѓ���������������̡�C�PL�BPQ�Ѓ����������������U���C�PL�EP�EPQ�JT�у�]� U���C�PL�EPQ��  �у�]� �U���C�PL�EPQ���   �у�]� ̡�C�PL�BXQ�Ѓ����������������U���C�PL�EP�EP�EPQ�J\�у�]� ������������U���4��CSV��HL�QW�ҋ�3ۉ}�;��x  �M�������C�E�EԋE�]Љ]؉]܉]�]��}̋Q�R0Ph]  �M��ҡ�C���   �BSSW���Ѕ���   ��C�QL�BW�Ћ���;���   ��    ��C���   �B(���ЍM�Qh�   ���u�����������   �M�;���   ��C���   ���   S��;�tm��C���   �ȋB<V�Ћ�C���   ���   �E�P�у�;�t��C�B@�HV�у���;��\����}��M�聹���M��I�����_^[��]� �}���C�B@�HW�ы�C���   ���   �M�Q�҃��M��9����M�����_^3�[��]� �����̡�C�PL�B`Q�Ѓ���������������̡�C�PL�BdQ�Ѓ����������������U���C�PL�EPQ�Jh�у�]� ���̡�C�PL��D  Q�Ѓ������������̡�C�PL�BlQ�Ѓ����������������U���C�PL�EPQ���   �у�]� �U��M��]�����U��M��U�@R��]��������������U��U�M��@R�UR��]����������U��U�M��@R�UR�UR�UR��]��U��U$�EV�Eh � h � h�� h�� R�Q�U R�UR�UR�U���A�$�5�C�vLRP���   Q�Ѓ�4^]�  ������̡�C�PL���   Q�Ѓ�������������U���C�PL�EP�EP�EPQ��   �у�]� ���������U���C�PL��H  ]�������������̡�C�PL��L  ��U���C�PL��P  ]��������������U���C�PL��T  ]��������������U���C�PL�EP�EP�EP�EP�EPQ���   �у�]� �U���C�PL�EP�EP�EPQ���   �у�]� ���������U���C�PL�EP�EP�EP�EPQ��   �у�]� �����U���C�HL���   ]��������������U���C�HL���   ]��������������U���C�HL���   ]�������������̡�C�HL��  ���C�HL��@  ��h4DPh^� � z  ���������������U��Vh4Dj\h^� ����y  ����t�@\��t
�MQV�Ѓ�^]� ������������U��� ��CV3��u��u�u�u�u��u��u􋈈   ���   W�ҋ}�E�;�t`;�t\��C�QLjP���   ���ЋM��U�Rh=���M�}���������C���   ���   �U�R�Ѓ��M��u��̴����_^��]Ë�C���   ���   �E�P�у��M��u�螴��_�   ^��]����U��� ��CV3��u��u�u�u�u��u��u􋈈   ���   W�ҋ}�E�;�t`;�t\��C�QLjP���   ���ЋM��U�Rh<���M�}��3�������C���   ���   �U�R�Ѓ��M��u��������_^��]Ë�C���   ���   �E�P�у��M��u��γ��_�   ^��]���̡�CV�񋈈   ���   V�҃��    ^��������������̡�CV��H�QV�ҡ�C�H$�QDV�҃���^�����������U���CV��H�QV�ҡ�C�H$�QDV�ҡ�C�U�H$�AdRV�Ѓ���^]� ��U���CV��H�QV�ҡ�C�H$�QDV�ҡ�C�U�H$�ARV�Ѓ���^]� ��U���CV��H�QV�ҡ�C�H$�QDV�ҡ�C�H$�U�ALVR�Ѓ���^]� �̡�CV��H$�QHV�ҡ�C�H�QV�҃�^�������������U���C�P$�EPQ�JL�у�]� ����U���C�P$�R]�����������������U���C�P$�Rl]����������������̡�C�P$�Bp����̡�C�P$�BQ�Ѓ����������������U���C�P$��VWQ�J�E�P�ы�C�u���B�HV�ы�C�B�HVW�ы�C�B�P�M�Q�҃�_��^��]� ���U���C�P$�EPQ�J�у�]� ����U���C�P$��VWQ�J �E�P�ы�C�u���B�HV�ы�C�B$�HDV�ы�C�B$�HLVW�ы�C�B$�PH�M�Q�ҡ�C�H�A�U�R�Ѓ� _��^��]� ���U���C�P$��VWQ�J$�E�P�ы�C�u���B�HV�ы�C�B$�HDV�ы�C�B$�HLVW�ы�C�B$�PH�M�Q�ҡ�C�H�A�U�R�Ѓ� _��^��]� ���U���,VW�E�P�o�����C�Q$�JP�E�P�ы�C�u���B�HV�ы�C�B�HVW�ы�C�B�P�M�Q�ҡ�C�H$�AH�U�R�Ћ�C�Q�J�E�P�у� _��^��]� �����̡�C�P$�B(Q��Yá�C�P$�BhQ��Y�U���C�P$�EPQ�J,�у�]� ����U���C�P$�EPQ�J0�у�]� ����U���C�P$�EPQ�J4�у�]� ����U���C�P$�EPQ�J8�у�]� ����U���C�UV��H$�ALVR�Ѓ���^]� ��������������U���C�H�QV�uV�ҡ�C�H$�QDV�ҡ�C�H$�U�ALVR�Ћ�C�E�Q$�J@PV�у���^]�U���C�UV��H$�A@RV�Ѓ���^]� ��������������U���C�P$�EPQ�J<�у�]� ����U���C�P$�EPQ�J<�у����@]� ���������������U���C�P$�EP�EPQ�JP�у�]� U���C�P$�EPQ�JT�у�]� ���̡�C�H$�QX�����U���C�H$�A\]�����������������U���C�P$�EP�EP�EPQ�J`�у�]� �����������̡�C�H(�������U���C�H(�AV�u�R�Ѓ��    ^]��������������U���C�P(�R]����������������̡�C�P(�B�����U���C�P(�R]�����������������U���C�P(�R]�����������������U���C�P(�R ]�����������������U���C�P(�E�RjP�EP��]� ��U���C�P(�E�R$P�EP�EP��]� ��C�P(�B(����̡�C�P(�B,����̡�C�P(�B0�����U���C�P(�R4]�����������������U���C�P(�RX]�����������������U���C�P(�R\]�����������������U���C�P(�R`]�����������������U���C�P(�Rd]�����������������U���C�P(�Rh]�����������������U���C�P(�Rx]�����������������U���C�P(�Rl]�����������������U���C�P(�Rt]�����������������U���C�P(�Rp]�����������������U�����C�E�    �E�    �P(�RhV�E�P���҅���   �E���uG��C�H�A�U�R�Ћ�C�Q�E�RP�M�Q�ҡ�C�H�A�U�R�Ѓ��   ^��]� ��C�Qh�h8  P���   �Ћ�C���E��Q(��u�B4j�����3�^��]� �M��Rj QP���҅�u�E�P�E����3�^��]� ��C�E��Q�M�j HP�EQ�JP�эU�R�tE�����   ^��]� �����U���C��V��H�A�U�R�Ѓ��M�Q������^��u��C�B�P�M�Q�҃�3���]� ��C�H$�E�I�U�RP�ы�C�B�P�M�Q�҃��   ��]� �U��Q��C�P(�RX�E�P�҅�u��]� �M3�8E�����   ��]� ���������U���C�P(�R8]�����������������U���C�P(�R<]�����������������U���C�P(�R@]�����������������U���C�P(�RD]�����������������U���C�P(�RH]�����������������U���C�P(�E�R|P�EP��]� ����U���C�P(�RL]�����������������U���C�E�P(�BT���$��]� ���U���C�E�P(�BPQ�$��]� ����̡�C�H(�Q�����U���C�H(�AV�u�R�Ѓ��    ^]��������������U���C�P(���   ]��������������U���C�H(�A]����������������̡�C�H,�Q,����̡�C�P,�B4�����U���C�H,�A0V�u�R�Ѓ��    ^]�������������̡�C�P,�B8�����U���C�P,�R<��VW�E�P�ҋu����C�H�QV�ҡ�C�H$�QDV�ҡ�C�H$�QLVW�ҡ�C�H$�AH�U�R�Ћ�C�Q�J�E�P�у�_��^��]� �������U���C�P,�E�R@��VWP�E�P�ҋu����C�H�QV�ҡ�C�H�QVW�ҡ�C�H�A�U�R�Ѓ�_��^��]� ��̡�C�H,�j j �҃��������������U���C�P,�EP�EPQ�J�у�]� U���C�H,�AV�u�R�Ѓ��    ^]�������������̡�C�P,�B����̡�C�P,�B����̡�C�P,�B����̡�C�P,�B ����̡�C�P,�B$����̡�C�P,�B(�����U���C�P,�R]�����������������U���C�P,�R��VW�E�P�ҋu����C�H�QV�ҡ�C�H$�QDV�ҡ�C�H$�QLVW�ҡ�C�H$�AH�U�R�Ћ�C�Q�J�E�P�у�_��^��]� �������U���C�H��D  ]��������������U���C�H��H  ]��������������U���C�H��L  ]��������������U���C�H�I]�����������������U���C�H�A]�����������������U���C�H�I]�����������������U���C�H�A]�����������������U���C�H�I]�����������������U���C�H���  ]��������������U���C�H�A]�����������������U���V�u�E�P���+�����C�Q$�J�E�P�у���u-��C�B$�PH�M�Q�ҡ�C�H�A�U�R�Ѓ�3�^��]Ë�C�Q�J�E�jP�у���u=�U�R��������u-��C�H$�AH�U�R�Ћ�C�Q�J�E�P�у�3�^��]Ë�C�B�HjV�у���u��C�B�HV�у����I�����C�Q$�JH�E�P�ы�C�B�P�M�Q�҃��   ^��]�����������U���C�H�A ]�����������������U���C�H�I(]�����������������U���C�H��  ]��������������U���C�H��   ]��������������U���C�H��  ]��������������U���C�H��  ]��������������U���C�H�A$��V�U�WR�Ћ�C�Q�u���BV�Ћ�C�Q$�BDV�Ћ�C�Q$�BLVW�Ћ�C�Q$�JH�E�P�ы�C�B�P�M�Q�҃�_��^��]������U���C�H���  ��V�U�WR�Ћ�C�Q�u���BV�Ћ�C�Q$�BDV�Ћ�C�Q$�BLVW�Ћ�C�Q$�JH�E�P�ы�C�B�P�M�Q�҃�_��^��]���U���C�H���  ]��������������U���<�<DSVW�E�    ��t�E�P�   �������/��C�Q�J�E�P�   �ы�C�B$�PD�M�Q�҃��}��C�H�u�QV�ҡ�C�H$�QDV�ҡ�C�H$�QLVW�҃���t)��C�H$�AH�U�R����Ћ�C�Q�J�E�P�у���t&��C�B$�PH�M�Q�ҡ�C�H�A�U�R�Ѓ�_��^[��]���U���C�H�U���  ��VWR�E�P�ы�C�u���B�HV�ы�C�B$�HDV�ы�C�B$�HLVW�ы�C�B$�PH�M�Q�ҡ�C�H�A�U�R�Ѓ� _��^��]����������������U��V�ujV�a�������^]���������̡�C�H���   ��U���C�H���   V�uV�҃��    ^]�������������U���C�P�]���C�P�B����̡�C�P���   ��U���C�P�R`]�����������������U���C�P�Rd]�����������������U���C�P�Rh]�����������������U���C�P�Rl]�����������������U���C�P�Rp]�����������������U���C�P�Rt]�����������������U���C�P���   ]��������������U���C�P�Rx]�����������������U���C�P���   ]��������������U���C�P�R|]�����������������U���C�P���   ]��������������U���C�P���   ]��������������U���C�P���   ]��������������U���C�P���   ]��������������U���C�P���   ]��������������U���C�P���   ]��������������U���C�P���   ]��������������U���C�P���   ]��������������U���C�P���   ]��������������U���C�P���   ]��������������U���C�P�EPQ��  �у�]� �U���C�P���   ]��������������U���C�P���   ]��������������U���C�P���   ]��������������U��E��t ��C�R P�B$Q�Ѓ���t	�   ]� 3�]� U���C�P �E�RLQ�MPQ�҃�]� U��E��u]� ��C�R P�B(Q�Ѓ��   ]� ������U���C�P�R]�����������������U���C�P�R]�����������������U���C�P�R]�����������������U���C�P�R]�����������������U���C�P�R]�����������������U���C�P�R]�����������������U���C�P�E�R\P�EP��]� ����U���C�E�P�B ���$��]� ���U���C�E�P�B$Q�$��]� �����U���C�E�P�B(���$��]� ���U���C�P�R,]�����������������U���C�P�R0]�����������������U���C�P�R4]�����������������U���C�P�R8]�����������������U���C�P�R<]�����������������U���C�P�R@]�����������������U���C�P�RD]�����������������U���C�P�RH]�����������������U���C�P�RL]�����������������U���C�P�RP]�����������������U���C�P���   ]��������������U���C�P�RT]�����������������U���C�P�EPQ��  �у�]� �U���C�P���   ]��������������U���C�P���   ]��������������U���C�P�RX]����������������̡�C�P���   ��U���C�P���   ]��������������U���C�P���   ]��������������U���C�P���   ]��������������U���C�P���   ]�������������̡�C�P���   ��U���C�P���   ]�������������̡�C�P���   ���C�P���   ���C�P���   ��U���C�H���   ]��������������U���C�H��   ]��������������U���C�H�U�E��VWRP���  �U�R�Ћ�C�Q�u���BV�Ћ�C�Q�BVW�Ћ�C�Q�J�E�P�у�_��^��]������������U���C�H���  ]��������������U���C�P(�} �R8����P��]� �U���C�P�BdS�]VW��j ���Ћ�C�Qh��p���   hc  V�Ћ�C���E��u�Q(�B4j�����_^3�[]� �Qj VP�Bh���Ћ�C�Q(�BHV���Ѕ�t ��C�Q(�E�R VP���҅�t�   �3��EP�0����_��^[]� ������U���C�U�� V��H$�IWR�E�P�ы�C���B�P�M�Q�ҡ�C�H�A�U�RW�Ћ�C�Q�J�E�P�у��U�R����������C�H�A�U�R�Ѓ�_��^��]� �����������h DPhD ��X  ���������������U��S�]W�;;�t_3�[]� V�s��u#��u9{u9yuP��uL9QuG^_�   []� �A��u��u9Qu��u'��u#9{�Յ�t��t;�u�C��tċI��t�;�t�^_3�[]� ���������U��EP�d������@]� �����������U��h DjhD �X  ����t
�@��t]��3�]��������Vh Dj\hD ����W  ����t�@\��tV�Ѓ���^�����Vh Dj`hD ���W  ����t�@`��tV�Ѓ�^�������U��Vh DjdhD ���yW  ����t�@d��t
�MQV�Ѓ�^]� ������������U��Vh DjhhD ���9W  ����t�@h��t
�MQV�Ѓ�^]� ������������Vh DjlhD ����V  ����t�@l��tV�Ѓ�^�������U��Vh Dh�   hD ����V  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh Dh�   hD ���vV  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh DjphD ���)V  ����t�@p��t�MQV�Ѓ�^]� �$D^]� ��U��Vh DjxhD ����U  ����t�@x��t
�MVQ�Ѓ���^]� ����������U��Vh DjxhD ���U  ����t�@|��t�MVQ�Ѓ�^]� 3�^]� �����U��Vh DjxhD ���iU  ����t�@|��t�MVQ�Ѓ����@^]� �   ^]� ������������̋���������������h DjhD �U  ����t	�@��t��3��������������U��V�u�> t+h DjhD ��T  ����t�@��tV�Ѓ��    ^]�������U��VW�}���t0h DjhD �T  ����t�@��t�MQWV�Ѓ�_^]� _3�^]� ����������U��Vh DjhD ���IT  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����U��Vh DjhD ���	T  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����Vh Dj hD ����S  ����t�@ ��tV�Ѓ�^�3�^���Vh Dj$hD ���S  ����t�@$��tV�Ѓ�^�3�^���U��Vh Dj(hD ���iS  ����t�@(��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vh Dj,hD ���S  ����t�@,��t�M�UQRV�Ѓ�^]� 3�^]� �U��Vh Dj(hD ����R  ����t�@0��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������Vh Dj4hD ���R  ����t�@4��tV�Ѓ�^�3�^���U��Vh Dj8hD ���YR  ����t"�@8��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���������U��Vh Dj<hD ���	R  ����t�@<��t
�MQV�Ѓ�^]� ������������Vh DjDhD ����Q  ����t�@D��tV�Ѓ�^�3�^���U��Vh DjHhD ���Q  ����t�M�PHQV�҃�^]� U��Vh DjLhD ���iQ  ����u^]� �M�PLQV�҃�^]� �����������U��Vh DjPhD ���)Q  ����u^]� �M�U�@PQRV�Ѓ�^]� �������Vh DjThD ����P  ����u^Ë@TV�Ѓ�^���������U��Vh DjXhD ���P  ����t�M�PXQV�҃�^]� U��Vh Dh�   hD ���P  ����u^]� �M�UQ�MR�UQ�MR���   QV�҃�^]� �����U��Vh Dh�   hD ���6P  ����u^]� �M�UQ�MR���   QV�҃�^]� �������������U��Vh Dh�   hD ����O  ����u^]� �M���   QV�҃�^]� �����U��Vh Dh�   hD ���O  ����u^]� �M���   QV�҃�^]� �����U��Vh Dh�   hD ���fO  ����u^]� �M���   QV�҃�^]� �����U��Vh Dh�   hD ���&O  ����t�M�UQ�MR���   QV�҃�^]� ��U���Vh Dh�   hD ��N  ����u��C�H�u�QV�҃���^��]ËM���   WQ�U�R�Ћ�C�Q�u���BV�Ћ�C�Q�BVW�Ћ�C�Q�J�E�P�у�_��^��]��U��Vh Dh�   hD ���VN  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh Dh�   hD ���N  ����t���   ��t�MQ����^]� 3�^]� �U��Vh Dh�   hD ����M  ����t���   ��t�MQ����^]� 3�^]� �U��Vh Dh�   hD ���M  ����t���   ��t�MQ����^]� 3�^]� �Vh Dh�   hD ���IM  ����t���   ��t��^��3�^����������������U��Vh Dh�   hD ���M  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh Dh�   hD ���L  ����t���   ��t�MQ����^]� ��������U��Vh Dh�   hD ���vL  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������Vh Dh�   hD ���)L  ����t���   ��t��^��3�^����������������VW��3����$    �h DjphD ��K  ����t�@p��t	VW�Ѓ���$D�8 tF��_��^�������U��SW��3�V��    h DjphD �K  ����t�@p��t	WS�Ѓ���$D�8 tqh DjphD �]K  ����t�@p��t�MWQ�Ѓ�����$Dh DjphD �+K  ����t�@p��t	WS�Ѓ���$DV���7�����tG�]����E^��t�8��~=h DjphD ��J  ����t�@p��t	WS�Ѓ���$D�8 u_�   []� _3�[]� ����������U��Vh Dj\hD ���J  ����t3�@\��t,V��h DjxhD �gJ  ����t�@x��t
�MVQ�Ѓ���^]� ��������U��Vh Dj\hD ���)J  ����t3�@\��t,V��h DjdhD �J  ����t�@d��t
�MQV�Ѓ���^]� ��������U���Vh Dj\hD ����I  ����tG�@\��t@V�ЋEh DjdhD �E��E�    �E�    �I  ����t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vh Dj\hD ���II  ����t\�@\��tUV��h DjdhD �'I  ����t�@d��t
�MQV�Ѓ�h DjhhD ��H  ����t�@h��t
�URV�Ѓ���^]� ���������������U��Vh Dj\hD ���H  ������   �@\��t~V��h DjdhD �H  ����t�@d��t
�MQV�Ѓ�h DjhhD �jH  ����t�@h��t
�URV�Ѓ�h DjhhD �AH  ����t�@h��t
�MQV�Ѓ���^]� ��U���Vh DjthD ���H  ����tQ�@t��tJ�MQ�U�VR�Ћu��P���?���h Dj`hD ��G  ����th�@`��ta�M�Q�Ѓ���^��]� h Dj\hD �G  �u����t4�@\��t-V��h DjdhD �xG  ����t�@d��th$DV�Ѓ���^��]� ������U���Vh Dh�   hD ���3G  ����tR���   ��tH�MQ�U�R���ЋuP���k���h Dj`hD ��F  ����t|�@`��tu�M�Q�Ѓ���^��]� h Dj\hD �E�    �E�    �E�    �F  �u����t3�@\��t,V��h DjdhD �F  ����t�@d��t
�U�RV�Ѓ���^��]� ��������������U���C���   �BXQ�Ѓ���u]� ��C�Q|�M�RQ�MQP�҃�]� ���U���C���   �BXQ�Ѓ���u]� ��C�Q|�M�R8Q�MQP�҃�]� ���U��EV��j ���C�Qj j P�B�ЉF����^]� ��̡�CVj ��H��Aj j R�Ѓ��F^����������������U��V��F��u^]� ��C�Q�MP�EP�Q�JP�у��F�   ^]� ���̡�C�H���   ��U���C�H���   V�u�R�Ѓ��    ^]����������̡�C�P���   Q�Ѓ�������������U���C�P�EPQ���   �у�]� ̡�C�H�������U���C�H�AV�u�R�Ѓ��    ^]��������������U���C�H�AV�u�R�Ѓ��    ^]��������������U���C�P��Vh�  Q���   �E�P�ы�C���   �Q8P�ҋ��C���   ��U�R�Ѓ���^��]��������������̡�C�P�BQ�Ѓ����������������U���C�P�EPQ�J\�у�]� ����U���C�P�EP�EP�EP�EP�EPQ���   �у�]� �U���C�P�EP�EP�EP�EPQ�JX�у�]� �������̡�C�P�B Q��Y�U���C�P�EP�EP�EP�EPQ���   �у�]� �����U���C�P�EP�EP�EPQ�J�у�]� ������������U���C�H��   ]��������������U���C�P�R$]�����������������U���C�P�EP�EP�EP�EPQ�J(�у�]� ��������U���C�P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ�J`�у�(]�$ ����U���C�P�EP�EP�EP�EPQ�J,�у�]� ��������U���CV��H�QWV�ҍx���C�H�QV�ҋ�C�Q�M�R4Q�MQ�MQWHPj j V�҃�(_^]� ���������������U���C�P�E P�EP�EP�EP�EP�EP�EPQ�J4�у� ]� ������������U���C�P�EP�EPQ�J@�у�]� U���C�P�EPQ�JD�у�]� ���̡�C�P�BLQ�Ѓ���������������̡�C�P�BLQ�Ѓ���������������̡�C�P�BPQ�Ѓ����������������U���C�P�EPQ�JT�у�]� ����U���C�P�EPQ�JT�у�]� ����U���C�P�EP�EPQ���   �у�]� �������������U���C�P�E���   ��VP�EPQ�M�Q�ҋu�    �F    ��C���   j P�BV�Ћ�C���   �
�E�P�у� ��^��]� ������̡�C�P�BhQ�Ѓ������������������3��Yp��A`�Ad�Ah�Ax�����A|   ����������������U��E��t�Ap��yd t�Ah]� 3��y|��]� ������̡�C�H�������U���C�H�AV�u�R�Ѓ��    ^]��������������U���C�P�E P�EP�EP�EP�EP�EP�EPQ�J�у� ]� ������������U���C�P�EPQ�J�у�]� ���̡�C�P�BQ��Y�U���C�P�EP�EPQ�J�у�]� U��VW���R���M�U�x@�EPQR���R���H ���_^]� �U��VW���R���M�U�xD�EPQR���nR���H ���_^]� �V���XR���xH u3�^�W���FR���΍xH�<R���H �_^�����U��V���%R���xL u3�^]� W���R���M�U�xL�EPQR����Q���H ���_^]� �������������U��V����Q���xP u���^]� W���Q���M�U�xP�EP�EQRP���Q���H ���_^]� ��������U��V���Q���xT u���^]� W���oQ���M�xT�EPQ���]Q���H ���_^]� U���S�]VW���t.�M��&������/Q���xL�E�P���!Q���H ��ҍM��`����}��tZ��C�H�A�U�R�Ћ�C�Q�J�E�WP�ы�C�B�P�M�Q�҃�����P���@@��t��C�QWP�B�Ѓ�_^[��]� ������U��VW���P���xH�EP���P���H ���_^]� ���������U��VW���dP���M�U�xD�EP�EQRP���JP���H ���_^]� �������������U��V���%P���xP u
�����^]� W���P���M�U�xP�EP�EQ�MR�UPQR����O���H ���_^]� ��������������U��V����O���xT u
�����^]� W���O���M�xT�EPQ���O���H ���_^]� ��������������U��V���uO���xX tW���gO���xX�EP���YO���H ���_^]� ������������U����MV3��E�PQ�u�u��u�u��u�u��h`  ����t.�E�;�t'��C�J�U�R�U�R�U�R�U�RP�AX�Ѓ�^��]�3�^��]������������̡�C�H��   ��U���C�H��$  V�u�R�Ѓ��    ^]�����������U���C�UV��H��(  VR�Ѓ���^]� �����������U���C�P�EQ��,  P�у�]� �U���C�P�EQ��,  P�у����@]� �����������̡�C�H��0  ���C�H��4  ��U��E��t�@�3���C�RP��8  Q�Ѓ�]� �����U���C�P�EPQ��<  �у�]� �U���C�P�EP�EP�EPQ��@  �у�]� ���������U���C�P�EP�EPQ��D  �у�]� �������������U���C�P�EPQ��H  �у�]� �U���C�P�E��L  ��VWPQ�M�Q�ҋu����C�H�QV�ҡ�C�H�QVW�ҡ�C�H�A�U�R�Ѓ�_��^��]� ��������������̡�C�P��T  Q�Ѓ������������̡�C�P��P  Q�Ѓ�������������U���C�P�EPQ��X  �у�]� ̡�C�H��\  ��U���C�H��`  V�u�R�Ѓ��    ^]�����������U���C�P�EP�EP�EP�EP�EPQ��d  �у�]� �U���C�P�EP�EP�EP�EP�EPQ��h  �у�]� �VW���O蔿����3��G �G$�G(�G,�G0�G4�G8�G<�G@�GD�GH�GL�GP�GT�GX�G\�_p��G`�Gd�Gh�Gx�����G|   ��_^����������������V��W�>��t7���/K���xP t$S���!K��j j �XPj�FP���K���H ���[�    �~` t��C�H�V`�AR�Ѓ��F`    _^������������U��SV��Fx��C�Q��   WV�^dSP�EP�~`W�у��F|����   �> ��   �; ��   �U�~pW�^hSR��^������u#���hX���C�H��0  h�   �҃��E�~P�������j j jW�N����F|��t��������F|_^[]� �F|_�Fx����^[]� �F|�����    ��C�Q��JP�у��    �F|_^[]� ���V��������3��^p��F`�Fd�Fh�Fx�����F|   ^�������U��QV��~d tg�E;Fxt_�N`W�>�M����{I���xP u����(S���hI���UR�XP�E�Pj�NQ���PI���H ���[�F|_��u�E�Fx�E��t�    �F`^��]� �M�Fx������t�3�^��]� ���������U��QVW�}�����\  ��C�H�QhV�҃�����Cu"�H��0  hX�h�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���t�3�9u�~�E���<� t��Q���Z  �EF;u�|�UR�M����_�   ^��]� �������������U��QVW�}����.\  ��C�H�QhV�҃�����Cu"�H��0  hX�h�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���tЋE��t�3�9u�~8��E�<� t'����C�QP�Bh�Ѓ���t�M��R���Y  F;u�|ʍEP�m
����_�   ^��]� �������������hX�h�   hPDh�   �7������t������3��������V��������N^��������������������U��VW�}�7��t�������N�ӻ��V������    _^]á�C�PD�BQ�Ѓ���������������̡�C�PD�BQ�Ѓ���������������̡�C�PD�BQ�Ѓ����������������U���C�PX��Q�
�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ���������U���C�PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U���C�PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U���C�PX��`VWQ�J�E�P�ы��E���   ���_^��]� �������������U���C�PX�EPQ�J�у�]� ����U���C�PX�EPQ�J�у�]� ����U���C�PX�EPQ�J�у�]� ����U���C�PX�EPQ�J�у�]� ����U���C�PX�EPQ�J$�у�]� ����U���C�PX�EPQ�J �у�]� ����U���C�PD�EP�EPQ�J�у�]� U���C�HD�U�j R�Ѓ�]�������U���C�H@�AV�u�R�Ѓ��    ^]��������������U���C�HD�	]��U���C�H@�AV�u�R�Ѓ��    ^]��������������U���C�HD�U�j R�Ѓ�]�������U���C�H@�AV�u�R�Ѓ��    ^]��������������U���C�U�HD�Rh'  �Ѓ�]����U���C�H@�AV�u�R�Ѓ��    ^]�������������̡�C�HD�j h�  �҃�����������U���C�H@�AV�u�R�Ѓ��    ^]�������������̡�C�HD�j h:  �҃�����������U���C�H@�AV�u�R�Ѓ��    ^]��������������U���3��E��E���C���   �R�E�Pj�����#E���]�̡�C�HD�j h�F �҃�����������U���C�H@�AV�u�R�Ѓ��    ^]�������������̡�C�HD�j h�_ �҃�����������U���C�H@�AV�u�R�Ѓ��    ^]��������������U��E����u��]� �E���C�E�    ���   �R�E�Pj������؋�]� ̡�C�PD�B$Q�Ѓ���������������̡�C�PD�B(Q�Ѓ���������������̡�C�PD�BQ�Ѓ���������������̡�C�PD�B(Q�Ѓ���������������̡�C�PD�BQ�Ѓ���������������̡�C�PD�B(Q�Ѓ���������������̡�C�PD�BQ�Ѓ���������������̡�C�PD�B(Q�Ѓ���������������̡�C�PD�BQ�Ѓ���������������̡�C�PD�B(Q�Ѓ���������������̡�C�PD�BQ�Ѓ���������������̡�C�PD�B(Q�Ѓ���������������̡�C�PD�BQ�Ѓ���������������̡�C�PD�B(Q�Ѓ���������������̡�C�PD�BQ�Ѓ���������������̡�C�PD�B(Q�Ѓ���������������̡�C�PD�BQ�Ѓ���������������̡�C�PD�B(Q�Ѓ���������������̡�C�PD�BQ�Ѓ���������������̡�C�H\�������U���C�H\�AV�u�R�Ѓ��    ^]�������������̡�C�P\�BQ�Ѓ���������������̡�C�P\�BQ�Ѓ����������������U���C�P\�EPQ�J�у�]� ����U���C�P\�EP�EPQ�J�у�]� U���C�P\�EPQ�J�у�]� ���̡�C�P\�BQ�Ѓ����������������U���C�P\�EPQ�J �у�]� ����U���C�P\�EP�EPQ�J$�у�]� U���C�P\�EP�EP�EPQ�J(�у�]� ������������U���C�P\�EPQ�J0�у�]� ����U���C�P\�EPQ�J@�у�]� ����U���C�P\�EPQ�JD�у�]� ����U���C�P\�EPQ�JH�у�]� ���̡�C�P\�B4Q�Ѓ����������������U���C�P\�EP�EPQ�J8�у�]� U���C�P\�EPQ�J<�у�]� ����U���SVW�}��j �ωu�������C�H\�QV�҃���S������3���~=��I ��C�H\�U�R�U��EP�A(VR�ЋM��Q���h����U�R���]���F;�|�_^[��]� ���������������U���VW�}�E��P�������}� ��   ��C�Q\�BV�Ѓ��M�Q�������E���t]S3ۅ�~H�I �UR���e����E�P���Z����E;E�!����C�Q\P�BV�ЋE@���E;E�~�C;]�|�[_�   ^��]� _�   ^��]� U��M�A8��   �IXV�AP�I@���I�AP�I(�AX�I ���I0���A@�I �A8�I(���IH������������Dz�u�؋��������^��]���W���A�IX�AP�I�A8�I�A�I@�AP�I@�U��A8�IX�]������IH�����I0�����e��	����ݝx����A�I(�U��A�I �U��AX�I �]��AP�I(�����IH�E����	���������I�������]��A8�I(�A@�I �����	�������I���E��e��I0�������]��E��e����]����e��ˋE��x������]������]��AH�I@�A0�IX�����]��AX�I�AH�I(�����]��A0�I(�A@�I�����]��AP�I0�AH�I8�����]��AH�I �AP�I�����]��A8�I�A0�I �   �����]��_^��]����̋�3ɉ�H�H�H�V��V�����FP����3����F�F^��3���A�A�A����A�`�
�@�b�	���B�a�������U����   ��UV���q�U�W3��<��M��}��'	  S�]����  ��؋���M�U��>���U�@�U���� �U��@�@�B�@�������@���@�   ���]��E��U�;���  �w�����  �w�������F�܍B��   �U������������ˋP��R�э����]��B���B�P���R���U����E������]��E��M��E������������]��E����E����E��E��]����E��]����E��]����]����U��E��U�����B���B���U������������]��E����E����������E������E��E��]����E��]����E��]��]��U���E��U��R�э����N�B���B�P���R���U������������]��E����E����������E������E��E��]����E��]����E��]����U��E��]�����B���B���U����E��������]��E����E����������E������E��E��U����E��]����E��U��E��U��T����E�ɋU�����������;���   �ߍ���+�������͋�@�������O�]��@���]��@���U������M������]��E��E����E������E����������E��E��U����E��]����E��U��E��E��U�u�������������������������[�[�E�����������������]  ��������������Dz���������E��+������������������M����M��E������������������[H���[P���[X�E����E���������zu������������zh�����CP���CX���CH���CX�������cH���[���[ �[(�C(�KP�C �KX���CX�K�C(�KH���CH�K �CP�K�����[0�[8�[@��   ������������z]�CX���CP�����cH�CH���CP�������[�[ �[(�C(�KP�C �KX���CX�K�C(�KH���CH�K �CP�K�����[0�[8�[@�]�CP���CX�����CH���CX�����cP���[0���[8�[@�C8�KX�C@�KP���CH�K@�C0�KX���C0�KP�C8�KH�����[�[ �[(��$���SQ������E��U�   �����}��M������3�3��u��u���|)�A�����B�4�u�0u��u�p��J�u�u�U�E;�}�Q���E���u��U��1���@���K�I�E    ��C0�H���CH�H��� �K �C�@�K8���@�KP���C(��C�@�K@���CX�H�D��@�����U���]�� �K��C0�H���@�KH��� �K �C�@�K8���@�KP��� �K(�C�C@�H���CX�H���U����n  �A�������@�E����E   �E�
���������ɋEH���׋��@�E�Ѝ��K��C0�H���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���CX�H�E������������������������������E����]��E��]����]�׋��@�E�Ѝ��K��C0�H���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���CX�H�E@������]������M������������������������]��E��]��E��]�׋��@�E�Ѝ��K��C0�H���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���CX�H���]������M������������������������]��E�E����]���E����]��E��M����@�E�Ѝ��K��C0�H���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���CX�H���]������M������������������������U��E��]��E��U������������������9M|��[��_��^���؋�]� ���������ʋE�����׋��@�E�Ѝ��K��C0�H���CH�H���]�� �K �C�@�K8���@�KP���]��C(��C�C@�H���CX�H�E@�E���]����E��������������������M����������]��E��E�;��T�����[������_��^��]� �����h0DPh_� ��  ���������������h0Djh_� �  ����uË@����U��V�u�> t/h0Djh_� �  ����t��U�M�@R�Ѓ��    ^]���U��Vh0Djh_� ���I  ����t�@��t�MQ����^]� 3�^]� �������U��Vh0Djh_� ���	  ����t�@��t�MQ����^]� 3�^]� �������U��Vh0Djh_� ����  ����t�@��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh0Djh_� ���y  ����t�@��t�MQ����^]� 3�^]� �������U��Vh0Dj h_� ���9  ����t�@ ��t�MQ����^]� 3�^]� �������U��Vh0Dj$h_� ����  ����t�@$��t�MQ����^]� 2�^]� �������Vh0Dj(h_� ���  ����t�@(��t��^��3�^������Vh0Dj,h_� ���  ����t�@,��t��^��3�^������U��Vh0Dj0h_� ���Y  ����t�@0��t�MQ����^]� 3�^]� �������U��Vh0Dj4h_� ���  ����t�@4��t�M�UQR����^]� ���^]� ��Vh0Dj8h_� ����  ����t�@8��t��^��3�^������U��Vh0Dj<h_� ���  ����t�@<��t�MQ����^]� ��������������U��Vh0Dj@h_� ���i  ����t�@@��t�MQ����^]� ��������������U��Vh0DjDh_� ���)  ����t�@D��t�MQ����^]� 3�^]� �������U��Vh0DjHh_� ����  ����t�@H��t�MQ����^]� ��������������Vh0DjLh_� ���  ����t�@L��t��^��3�^������Vh0DjPh_� ���|  ����t�@P��t��^��3�^������Vh0DjTh_� ���L  ����t�@T��t��^��^��������Vh0DjXh_� ���  ����t�@X��t��^��^��������Vh0Dj\h_� ����  ����t�@\��t��^��^��������U��Vh0Dj`h_� ���  ����t�@`��t�M�UQR����^]� 3�^]� ���U��Vh0Djdh_� ���y  ����t�@d��t�M�UQR����^]� 3�^]� ���U��Vh0Djhh_� ���9  ����t�@h��t�M�UQ�MR�UQ�MRQ����^]� ��������������U��Vh0Djlh_� ����  ����t�@l��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh0Djph_� ���  ����t�@p��t�M�UQR����^]� 3�^]� ���U��Vh0Djth_� ���Y  ����t�@t��t�M�UQR����^]� 3�^]� ���U��Vh0Djxh_� ���  ����t�@x��t�M�UQR����^]� 3�^]� ���U��Vh0Dj|h_� ����  ����t�@|��t�MQ����^]� 3�^]� �������U��Vh0Dh�   h_� ���  ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh0Dh�   h_� ���F  ����t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh0Dh�   h_� ����  ����t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh0Dh�   h_� ���  ����t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U���|��A���U����U����U���  S�V�E��EW�����������   ���������U�r�z�
�R;��4v���4��I�$ȍ��F�R�a���F�a�uB�!�]��B�a�U��B�a�U������������]��E����E����������E��������E��G��$ȍ��]��B�a�U��B�a�U������������]��E����E����������E��������E��������M�������_�U�^��[�U����U���������������������M  ��������������D�Ez���P�P���]� �������E�����E����X�M��X��]� ����U���@����A���E�    �����]����]��]�����������]����]��]����   �	S�]VW�M��E����������t[��%�����E�M�����@��P�}����F�@��R�M��k����~���Q�M��Y����v;�t�v��P�M��C����M����M��M�u��}� _^[tV�E؋E�E����E��E����E��E����8�������������X���X��� ���`���`�E����X�X��]� ��E����������P���P�E����X�X��]� �����������̋Q3���|�	��t��~�    t@��Ju��3�����������U��QV�u��;�}�	���    u@��;�|����^]� +�@^]� �����������U��VW�}��x+�1��t%�Q3���~�΍I �1�������;�t@��;�|���_^]� �Q3���~!V�1�d$ ���   @u	�����t@��Ju�^�����̋QV3���~�	�d$ ����ШtF��Ju��^�����������U��Q3�9A~��I ��$������@;A|�Q��~YSVW�   3ۋ���x5��%����E���;�}$�I �������%���;E�u�
   �F;q|ߋQG�G���;�|�_^[��]�����������U��	����%�����E��   @t������A��wg�$�Xb�E�M� �������]� ��M��P�E�]� �H�U�
�@�M�]� �P�M��P�E�]� �H�U�
� �M�]� ���abb/bCb����U����S��V�����W�   @t���������];�t�����u�};�tK�����tC��}�����t�������t�Ӄ��t��_%   ��^�[]� �%   ���   @�_^[]� ����V��V�����FP����3����F�F^��U��SV��WV�r����^S�i����E3����~�~;�t_��C�Q���   h����jIP�у��;�t9�}��t;��C�B���   h����    jNQ�҃����uV�������_^3�[]� �E�~_�F^�   []� ����������U��V��WV������FP�����}���F    �F    ����   �? ��   �G����   ��C�Q���  h����jlP�у����t>� t@�G��t9��C�Jh����    ���  jqR�Ѓ��F��u���v���_3�^]� �O��N�G�F��    ���t��t��tQPR�SZ  ���F��t�VP��RP�GP�  ��_�   ^]� ��������U��SV��WV�����~W����3����F�F9E�  �];���   ��C�Qh����    h�   P���  �Ѓ����t@�} tN�]��tD��C�Q���  h����    h�   P�у����u���n���_^3�[]� �^�]�0�]�F   ��C�B���  h��h�   j�у����t���^��t��    ��t�UQRP�Y  ���E��t!�N�?�W�QWP�R  ��_^�   []� ��_^�   []� ���U��Q�A�E� ��~JS�]V�1W����$    ����������;�u�   @u�����u3��	�   ����U���Ou�_^[�E��Ћ�]� �����������U��S�]V��3�W�~���F�F�CV;C��   �����W�����3��F�F��C�Q���   h��jIj�Ѓ������   ��C�Q���   h��jNj�Ѓ����uV������_��^[]� ��F   �F   ����K�H�C��B�_��^�   []� �@���W�:���3��F�F��C�B���   h��jIj�у����t[��C�B���   h��jNj�у�����\�����F   �F   ����S�Q��K�H��C�B��   _��^[]� �����������U��3�V���F�F�F�EP������^]� �������������U��EVP��������^]� ����������U��U��t�M��t�E��tPRQ�V  ��]�����������̋�3ɉH��H�@   �������������U��ыM��tK�E��t��C���   P�B@��]� �E��t��C���   P�BD��]� ��C���   R�PD��]� �����U���C�P@�Rd]�����������������U���C�P@�Rh]�����������������U���C�P@�Rl]�����������������U���C�P@�Rp]�����������������U���C���   ���   ]�����������U���C���   ���   ]����������̡�C�P@�Bt����̡�C�P@�Bx�����U���C�P@�R|]����������������̡�C�P@���   ���C���   �Bt��U���C�P@���   ]�������������̡�C�P@���   ��U���C�P@���   ]��������������U���C�P@���   ]��������������U���C�P@���   ]��������������U���C�P@���   ]��������������U���CV��H@�QV�ҋM����t��#�����C�Q@P�BV�Ѓ�^]� �̡�C�PH���   Q�Ѓ�������������U���C�P@�EPQ�JL�у�]� ���̡�C�P@�BHQ�Ѓ����������������U���C�P@�EP�EP�EPQ�J�у�]� ������������U���C�P@�EPQ�J�у�]� ����U���C�P@�EP�EPQ�J�у�]� U���C�P@�EPQ�J �у�]� ����U���C���   �R]��������������U���C���   �R]��������������U���C���   �R ]��������������U���C���   ���   ]�����������U���C���   ��D  ]�����������U���C�E���   �E ���   P�E���$P�EP�EP�EP��]� ���������U���C���   ���   ]����������̡�C���   �B$���C�H@�Q0�����U���C�H@�A4j�URj �Ѓ�]����U���C�H@�A4j�URh   @�Ѓ�]�U���C�H@�U�E�I4RPj �у�]�̡�C�H|�������U��V�u���t��C�Q|P�B�Ѓ��    ^]��������̡�C�H|�Q �����U��V�u���t��C�Q|P�B(�Ѓ��    ^]��������̡�C�H@�Q0�����U��V�u���t��C�Q@P�B�Ѓ��    ^]���������U���C�H@���   ]��������������U��V�u���t��C�Q@P�B�Ѓ��    ^]��������̡�C�PH���   Q�Ѓ�������������U���C�PH�EPQ��d  �у�]� �U���C�H �IH]�����������������U��}qF uHV�u��t?��C���   �BDW�}W���Ћ�C�Q@�B,W�Ћ�C�Q�M�Rp��VQ����_^]����������̡�C�P@�BT�����U���C�P@�RX]�����������������U���C�P@�R\]����������������̡�C�P@�B`�����U���C�H��T  ]��������������U���C�H@�U�A,SVWR�Ћ�C�Q@�J,���EP�ы�C�Z��h��hE  �΋��g��Ph��hE  ����f��P��T  �Ѓ�_^[]����U��E�M�UP��P�EjP��(����]��������������̸   �����������U��V�u��t���u6�EjP��(������u3�^]Ë��)����t���t��U3�;P��I#�^]�������h4DPh^� �������������������U��Vh4Djh^� ���y�������t�@��t�M�UQRV�Ѓ�^]� 3�^]� �Vh4Djh^� ���<�������t�@��tV�Ѓ�^�3�^���U��Vh4Djh^� ���	�������t�@��t�M�UQRV�Ѓ�^]� ���^]� U���  Vh4Djh^� �����������t/�@��t(�MWQ��x���VR�Ћ��E���b   ���_^��]� �u���3����N`�+������   � �����   ������ݞ�  ��^��]� ����U��Vh4Djh^� ���9�������t�@��t�M�UQRV�Ѓ�^]� ��������U��Vh4Djh^� �����������t�@��t�M�UQ�MRQV�Ѓ�^]� ����U��Vh4Dj h^� ����������t�@ ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vh4Dj$h^� ���i�������t�@$��t�MQV�Ѓ�^]� 3�^]� �����U��Vh4Dj(h^� ���)�������t�@(��t�M�UQ�MR�UQRV�Ѓ�^]� U��QVh4Dj,h^� �����������t �@,�E���t�E�MPQV�U���^��]� ��^��]� ��������U��Vh4Dj0h^� ����������t#�@0��t�E�M�U���$QRV�Ѓ�^]� 3�^]� ��������Vh4Dj4h^� ���L�������t�@4��tV�Ѓ�^�3�^���Vh4Dj8h^� ����������t�@8��tV�Ѓ�^�������U���`Vh4DjDh^� �����������t(�@D��t!W�M�VQ�Ћ��E���   ���_^��]� �u���]�����^��]� ����U��Vh4DjHh^� ����������t�@H��t
�MQV�Ѓ�^]� ������������U��Vh4DjLh^� ���I�������t�@L��t�MQV�Ѓ�^]� ���^]� ����U��Vh4DjPh^� ���	�������t�@P��t
�MQV�Ѓ�^]� ������������U��Vh4DjTh^� �����������t�@T��t
�MQV�Ѓ�^]� ������������U��Vh4DjXh^� ����������t.�@X��t'�M �UQ�MR�UQ�MR�UQ�MRQV�Ѓ� ^]� 3�^]� �������������Vh4Dj`h^� ���,�������t�@`��tV�Ѓ�^�3�^���U��Vh4Djdh^� �����������t�@d��t�MQV�Ѓ�^]� 3�^]� �����U���Vh4Djhh^� ����������t1�@h��t*�MQ�U�VR�Ћu��P�������M��ǡ����^��]� �u��脡����^��]� �����������Vh4Djph^� ���L�������t�@p��tV�Ѓ�^Ã��^��Vh4Djlh^� ����������t�@l��tV�Ѓ�^Ã��^��Vh4Djth^� �����������t�@t��tV�Ѓ�^�3�^���U��Vh4Djxh^� ����������t�@x��t
�MQV�Ѓ�^]� ������������Vh4Dj|h^� ���|�������t�@|��tV�Ѓ�^�������Vh4Dh�   h^� ���I�������t���   ��tV�Ѓ�^�U��Vh4Dh�   h^� ����������t���   ��t�MQV�Ѓ�^]� ���^]� ��������������U��Vh4Dh�   h^� �����������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U���Vh4Dh�   h^� ���s�������tU���   ��tKW�M�VQ�Ћ�C�u���B�HV�ы�C�B�HVW�ы�C�B�P�M�Q�҃�_��^��]� ��C�H�u�QV�҃���^��]� ����������Vh4Dh�   h^� �����������t���   ��tV�Ѓ�^Ã��^������������U��Vh4Dh�   h^� ����������t���   ��t
�MQV�Ѓ�^]� ������U��Vh4Dh�   h^� ���V�������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh4Dh�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������Vh4Dh�   h^� ����������t���   ��tV�Ѓ�^�3�^�������������U��Vh4Dh�   h^� ���v�������t%���   ��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���U��Vh4Dh�   h^� ���&�������t���   ��t�M�UQRV�Ѓ�^]� ���^]� ����������U��Vh4Dh�   h^� �����������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh4Dh�   h^� ����������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh4Dh�   h^� ���6�������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh4Dh�   h^� �����������t���   ��t�MQV�Ѓ�^]� ���^]� ��������������Vh4Dh�   h^� ����������t���   ��tV�Ѓ�^�3�^�������������Vh4Dh�   h^� ���Y�������t���   ��tV�Ѓ�^�3�^�������������Vh4Dh�   h^� ����������t���   ��tV�Ѓ�^�3�^�������������Vh4Dh�   h^� �����������t���   ��tV�Ѓ�^�3�^�������������U��Vh4Dh�   h^� ����������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������Vh4Dh�   h^� ���I�������t���   ��tV�Ѓ�^�3�^�������������U���Vh4Dh�   h^� ����������tF���   ��t<�MQ�U�VR�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ��U��Vh4Dh�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� ��Vh4Dh�   h^� ���I�������t���   ��tV�Ѓ�^�3�^�������������U���Vh4Dh�   h^� ����������tF���   ��t<�MQ�U�VR�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ��U��Vh4Dh�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� ��Vh4Dh�   h^� ���I�������t���   ��tV�Ѓ�^�3�^�������������U��Vh4Dh�   h^� ����������t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��QVh4Dh�   h^� ����������t#���   �E���t�E�MPQV�U���^��]� ��^��]� ��U��Vh4Dh�   h^� ���f�������t!���   ��t�E�M�U���$QRV�Ѓ�^]� ���������U��Vh4Dh�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh4Dh�   h^� �����������t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh4Dh   h^� ���v�������t��   ��t�MQV�Ѓ�^]� 3�^]� ���������������Vh4Dh  h^� ���)�������t��  ��tV�Ѓ�^�3�^�������������U���Vh4Dh  h^� �����������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U���Vh4Dh  h^� ���c�������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U���Vh4Dh  h^� �����������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U��Vh4Dh  h^� ���f�������t��  ��t
�MQV�Ѓ�^]� ������U��Vh4Dh  h^� ���&�������t��  ��t
�MQV�Ѓ�^]� ������U��Vh4Dh  h^� �����������t��  ��t
�MQV�Ѓ�^]� ������Vh4Dh   h^� ����������t��   ��tV�Ѓ�^�3�^�������������U��Vh4Dh$  h^� ���f�������t��$  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh4Dh(  h^� ����������t!��(  ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh4Dh,  h^� �����������t��,  ��t�M�UQ�MRQV�Ѓ�^]� ��������������Vh4Dh0  h^� ���y�������t��0  ��tV�Ѓ�^�3�^�������������U��Vh4Dh4  h^� ���6�������t��4  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh4Dh8  h^� �����������t��8  ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh4Dh<  h^� ����������t��<  ��t�M�UQ�MRQV�Ѓ�^]� ��������������U��Vh4Dh@  h^� ���F�������t��@  ��t�M�UQ�MRQV�Ѓ�^]� ��������������Vh4DhD  h^� �����������t��D  ��tV�Ѓ�^�3�^�������������U��Vh4DhH  h^� ����������t��H  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh4DhL  h^� ���f�������t��L  ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh4DhP  h^� ����������t!��P  ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��QVh4DhT  h^� �����������t'��T  �E���t�E�M�UPQRV�U���^��]� ��^��]� ��������������U��Vh4DhX  h^� ���f�������t%��X  ��t�E�M�U���$Q�MRQV�Ѓ�^]� �����U��Vh4Dj<h^� ����������t�@<��t�M�UQRV�Ѓ�^]� ��������U��Vh4Dj@h^� �����������t�@@��t�MQV�Ѓ�^]� 3�^]� �����h8DPh�� �������������������h8Djh�� ��������uË@����U��V�u�> t/h8Djh�� �S�������t��U�M�@R�Ѓ��    ^]���U��Vh8Djh�� ����������t �@��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh8Djh�� �����������t�@��t�M�UQR����^]� ����������U��Vh8Djh�� ����������t�@��t�M�UQR����^]� ����������U��Vh8Djh�� ���I�������t(�@��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��Vh8Dj h�� �����������t$�@ ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �������U��Vh8Dj$h�� ����������t �@$��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh8Dj(h�� ���Y�������t �@(��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh8Dj,h�� ���	�������t0�@,��t)�M$�E�UQ�M���\$�E�$R�UQR����^]�  3�^]�  �����������U��Vh8Dj0h�� ����������t$�@0��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �������U��Vh8Dj4h�� ���Y�������t5�@4��t.�M(�E �UQ�M���$R�UQ�MR�UQ�MRQ����^]�$ 3�^]�$ ������U��QVh8Dj8h�� �����������t�@8�E���t�E�MPQ���U�^��]� ��^��]� ����������U��Vh8Dj<h�� ����������t�@<��t�M�UQR����^]� ����������U��Vh8Dj@h�� ���i�������t�@@��t�M�UQR����^]� 3�^]� ���U��Vh8DjHh�� ���)�������t�@H��t�M�UQR����^]� 3�^]� ���U��Vh8DjDh�� �����������t�@D��t�M�UQR����^]� 3�^]� ���U��QVh8DjLh�� ����������t#�@L�E���t�E�EP�����$�U�^��]� ��^��]� �����U��Vh8DjPh�� ���Y�������t�@P��t�M�UQR����^]� 3�^]� ���U��Vh8DjTh�� ����������t �@T��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh8DjXh�� �����������t(�@X��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��Vh8Dj\h�� ���y�������t(�@\��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��V��~ Wu h8Djh�� �"�������t�@�ЉF�~��t6h8Djh�� ���������t�@��t�M�UVQ�MRQ����_^]� _3�^]� ��������������U��V��W�~��t+h8Djh�� ��������t�@��t�M�UQR���Ѓ~ t1h8Djh�� �p�������t�N�U�M�@R�Ѓ��F    _^]� ����������U��V��~ u h8Djh�� �#�������t�@�ЉF�v��t+h8Djh�� ���������t�@��t�M�UQR����^]� �������������U��V�q��t@h8Djh�� ��������t(�@��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ��������������U��V�q��t<h8Dj h�� �T�������t$�@ ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� ��U��SV��~ Wu h8Djh�� ��������t�@�ЉF�}�]�M�UWSQR���  ��t;�v��t4h8Dj$h�� ��������t�@$��t�M�UWSQR����_^[]� _^3�[]� ���U��V�q��t8h8Dj(h�� �t�������t �@(��t�M�UQ�MR�UQR����^]� 3�^]� ������U��V�q��tHh8Dj,h�� �$�������t0�@,��t)�M$�E�UQ�M���\$�E�$R�UQR����^]�  3�^]�  ������U��V�q��t<h8Dj0h�� ���������t$�@0��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� ��U��EHu�E�M�DD�@D�   ]� �������������U��EHV����   �$�$��   ^]áHD@�HD��uT�EP�7�����=�.  }�����^]Ëu��t�h�jmhPDj��������t ���d���<D��tV���\h���   ^]��<D    �   ^]ËM�UQR�5����������H^]�^]������HDu.�����>����<D��t���d��V�׵�����<D    �   ^]Ã��^]�@�ٔ��8��������hLDPh�f �0������������������U��hLDjh�f ��������t
�@��t]�����]�������U��VhLDjh�f �����������tC�~ t=�E8�M4�U0P�E,Q�M(RPQ���U��R�zc���E�NP�у�4�M���c����^]ÍM�c�����^]��U��hLDjh�f �l�������t
�@��t]��3�]��������U��hLDjh�f �<�������t�x t�P]��3�]������V��FW��u�~��N�<��u�< ��u_3�^á�C�H�F��  h@�j8��    RP�у���tщ~�F_�   ^���U��V��F;Fu������u^]� �N�V�E���   F^]� �����������U��S�]V��F;�~ ��x�F�M��^�   []� ^3�[]� }jW�F9FuK��u�~��N�<��u�< ��tA��C�B�V��  h@�j8��    QR�Ѓ���t�F�~�N�V��    �F9^|�_�F;Fu���������u����N�V�E���   F^[]� ��U��V��FW�};�~����y3�;Fu�m�����u_^]� �F;�~�N�T����H�;��F�M���F_�   ^]� ����U��E��x2�Q;�}+J�Q;�}V��    �Q�t���@�2;A|�^�   ]� 3�]� ��������������U��Q3�V��~�I�u91t@��;�|���^]� ���������V��W�~W����3����_�F�F^�����A    ��������̋Q�B���x;�}�QV�4���tP�1�����^�3�����������̍Q3��Q�Q�A�Q�A������������W���O�G;�t#��tV�q��t�~ u3���j�ҋ΅�u�^�G�G�G�G    �G�G    _�����U��A��3�V;�t��t�M��B;�t�@��t
�x t��u�3�^]� ����������U��Q�E�P�Q�P�Q�B�A]� �U��E�Q�P�Q�P�Q�B�A]� ̋Q��3�;�t�ʅ�t�I@��t
�y t��u�������������U��E�P�Q�H�A�@�H]� ����U��E�P�Q�H�A�A�H]� ���̋Q��t!�A��t�B�A�Q�P�A    �A    ��������V��W�~W�������3����_�F�F^��������������U���SV�uW���^S�}�趬��3���F�F�O�N�W���V�E9G~|��I �O���F�U�9FuL��u�~��~��t���< ��tY��C�H���  h@�j8��    RP�у���t0�~�}���V��M����E�F@�E;G|�_^�   [��]� _^3�[��]� U��V�u��x'�A;�} �U��x;�};�t�A��W�<��<���_^]� ���������U��EV�u;�}N��x,�Q;�}%��x!;�};�t�QW�<�P������tVW����_^]� ������������U��V�q3�W��~�Q�}9:t@��;�|����Ѕ�x);�}%N�q;�}�A�t���B�0;Q|�_�   ^]� _3�^]� ������U����E�Qj�E��ARP�M��E����[�����]� �����U����Q�Ej�E��A�MRPQ�M��E����w�����]� ̋A��;�t?W3�;�t7V�H;�t	9yt���3��P;�t;�t�J�H�P�Q�x�x��;�u�^_������̋Q�8���t!�A��t�B�A�Q�P�A    �A    �̋�� ���@8��HV3��q�q�P�r�r�8��p�p�p�P�H^������V������r����F3��F8�;�t�N;�t�H�F�N�H�V�V�F�F8�;�t�N;�t�H�F�N�H�V�V^�U��E�UP�AR�Ѓ�]� ���������U��V��N3��8�;�t�F;�t�A�F�N�H�V�V�Et	V�v�������^]� ������������U��V��W�~W����
���3����E��F�Ft	V�1�����_��^]� ������U��V��������Et	V�	�������^]� ���������������U���C�PH�EPQ���  �у�]� �U���C�P�B4VW�}j��h�  ���ЋMWQ���T  _^]� ��������������U��V���PXW�ҋ}P���|�����Et�_�   ^]� �M�UPWQR���A  _^]� �����������U��S�]VW��j ���z���8�  �}uI�~ uC��C�P���   j h�  ���Ѕ�u��C�QP���   h�  ���Ѕ�t	_^3�[]� �M�U�EQ�MRPSWQ����  _^[]� ��������U��EP�A    �]W����]� �����̸   �A� ������A   � ������U���@S�]VW����`��u�G   �y  ����   �M3�V�y���8�  u4�]N��P�w��V����C�P�M�B4��jh�  ��_^�C�[��]� �MV�Uy���8�  u�E�M��RPQ����_^�   [��]� �MV�%y���8�  t�MV�y���8��  ��C�P�M�B4jh�  �Љw�  ����  �E�H��BXj	��P����3��؃��u�;�t��C�QH���  VS�Ѓ��E��M�;O�b  9w�Y  ��C�B�M���   Vh�  �҅�u!��C�P�M���   Vh�  �Ѕ��  ��C�Q�M�B4Vh�  ��;�t
V���������E��G��C���   ���   �Ћ]�E�;���   ;���   S�T���M���jQ�ˉu��uĉuȉủuЉu؉u��B:���U�E��ˉu��u�u�U�E��]��E�   �\I����tHtHt�u���E�   ��E�   ��E�   �����M�;�t�M����BX�M�Q����P�_����M܃�;�t�M���M��8	���M��0	���M��hU���]�U�E�MRSPQ���  _^[��]� ��C���   ���   �E�P�у�_^�   [��]� ��������������̸   � ��������� ������������̃��� ����������� �������������U���C�H�QV�uV�҃���^]� ̸   � ��������3�� ����������̸   @� ��������3��  ����������̸   � ��������U��W�}��u3�_]� ��U�@@VR�Ћ���u^_]� ��C�Q0�F�M���   PQW�ҋF��^_]� U���C�H0�U�AR�Ѓ���t
��ȋj��]� �������3�� ��������������������������̸   � ��������3�� �����������3�� �����������U��E� ����]� �������������̸   � ��������U��E� ����]� ��������������3�� �����������U���C�H���  ]��������������U���C�H���  ]��������������U���C�P�EP�EP�EP�EPQ���   �у�]� �����U���C�E�P�EP�E���\$�E�$PQ���   �у�]� �������������U���C�P�EP�EP�EPQ���   �у�]� ��������̡�C�P���   Q�Ѓ�������������U���C�P�EP�EP�EPQ���   �у�]� ���������U���C�P�EP�EPQ���   �у�]� �������������U���C�H�U�ApR�Ѓ�]� �����U���C�P�EP�EPQ���  �у�]� �������������U���C�P�EP�EPQ���  �у�]� �������������U���C�P�EP�EPQ���  �у�]� �������������U���C�P�EP�EPQ���  �у�]� �������������U����   V�u��u3�^��]�Wh�   ��0���j P�4  ��R���E�P���ҡ�C�P�B<�M��Ћ}��t0j �M�QW��������u��C�B�P�M�Q�҃�_3�^��]ËE�M�Uh�   ��p�����0���P��t����MQWj	��P�����0���ǅ4����� �E�0��E�P��E����E��� �E�`� �E��� �E��� ǅx����� ǅ|��� ��E�`��E����E�P� �E�p��E����E���E�@� �E����E����E�@��Eİ� ������C���B�P�M�Q�҃�_��^��]����������U���   SV�u(3ۉ]���u��C�H�A�UR�Ѓ�^3�[��]Ë�C�Q�B<W�M3��Ѕ��N  �l����E�����   �MQ�M��O����C�B�P�M�Q�ҡ�C�H�AWj��U�hl�R�Ѓ��M�Q�M��kO���u�Wj��U�R�E�P��\���Q�_?��a����P��x���R�^S����P�E�P�QS����P��膃���E���t�E� �� t�M�����O����t��x�������vO����t��\�������cO����t�M̃���SO����t��C�Q�J�E�P����у���t�M��)O���}� t"�U(�E$�M�R�UP�EQ�MRPQ����������U�R�8�������E$�M�UVP�Ej QRP�����������C�Q�J�EP�у���_^[��]���������U��E�M�UP�EQ�Mj RPQ������]�������������̋�`L����������̋�`����������̋�` ����������̋�`����������̋�`$����������̋�`4����������̋�`D����������̋�`T����������̋�`����������̋�`(����������̋�`8����������̋�`H���� 2�2���2<��2u��2���2�2
��2��� 2\��$2��Ë�U�������} t�!  ��]��̃��$�m$  �   ��ÍT$�$  R��<$�D$tQf�<$t��#  �   �u���=TD �C$  �   ��1�@$  �  �u,��� u%�|$ u���#  �"��� u�|$ u�%   �t����-��   �=TD ��#  �   ��1��"  ZË�Q����$  YË�U��V��������EtV轝��Y��^]� ����̃=tb t-U�������$�,$�Ã=tb t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$������̋T$�L$��ti3��D$��u���   r�=tb t�'  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$�������U��WV�u�M�}�����;�v;���  ���   r�=tb tWV����;�^_u�.'  ��   u������r)��$�Я�Ǻ   ��r����$���$����$�d���� �D�#ъ��F�G�F���G������r���$�Я�I #ъ��F���G������r���$�Я�#ъ���������r���$�Я�I ǯ���������������D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�Я��������E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�l������$���I �Ǻ   ��r��+��$�p��$�l������̰�F#шG��������r�����$�l��I �F#шG�F���G������r�����$�l���F#шG�F�G�F���G�������V�������$�l��I  �(�0�8�@�H�P�c��D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�l���|��������E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_��jh "�s4  �E��uz�.4  ��u3��8  �R(  ��u�34  ����3  ���xb�3  �\D�H-  ��y��$  ���F2  ��x ��/  ��xj �
+  Y��u�XD��   �T/  ��3�;�u[9=XD~��XD�}�9=�Ju�,  9}u�$/  �$  �3  �E������   �   3�9}u�=42�t�n$  ��j��uY�-$  h  j�6)  YY��;�����V�542�5�J� ��Ѕ�tWV�f$  YY����N��V��  Y�������uW�&  Y3�@�c3  � jh@"�3  ����]3�@�E��u9XD��   �e� ;�t��u.�����tWVS�ЉE�}� ��   WVS�C����E����   WVS�_����E��u$��u WPS�K���Wj S���������tWj S�Ѕ�t��u&WVS�������u!E�}� t�����tWVS�ЉE��E������E���E��	PQ�s5  YYËe��E�����3��k2  Ë�U��}u�n5  �u�M�U�����Y]� ��U��S�]���woVW�=�K u�d   j�  h�   �T(  YY��t���3�@Pj �5�K������u&j^9 LtS�.6  Y��u����5  �0��5  �0��_^�S�6  Y�5  �    3�[]Ë�U��} t-�uj �5�K����uV�~5  ����P�.5  Y�^]����̃=La ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU��5  ��=La t2���\$�D$%�  =�  u�<$f�$f��f���d$u�5  ���$�"  �   ��ÍT$��  R��<$tmf�<$t�  =  �?s+��������������=TD ��  �   ��1��  w:�D$��%�� D$u)��   ����-�t�����B  ���� u�|$ u����-��   �=TD ��  �   ��1�  Z����������̃=La ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�	:  ��=La t2���\$�D$%�  =�  u�<$f�$f��f���d$u�9  ���$��  �   ��ÍT$�}  R��<$tmf�<$t�9  =  �?s-����������������=TD ��  �   ��1�  w8�D$��%�� D$u'��   ���t���������  ���� u�|$ u����-��   �=TD �:  �   ��1�C  Z����������̃=La ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�>  ��=La t2���\$�D$%�  =�  u�<$f�$f��f���d$u��=  ���$�  �   ��ÍT$�-  R��<$tPf�<$t�-H�������z�=TD �\  �   ��1�Y  �-J���������z��������  ���� u�|$ u����-��   �=TD �  �   ��1�  Z�������̃=La ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�>  ��=La t2���\$�D$%�  =�  u�<$f�$f��f���d$u�E>  ���$�R  �   ��ÍT$��  R��<$tPf�<$t�-H�������z�=TD �,  �   ��1�)  �-J���������z��������  ���� u�|$ u����-��   �=TD ��  �   ��1��  Z�������̃=La �B  ���\$�D$%�  =�  u�<$f�$f��f���d$��A  � �~D$f(��f(�f(�fs�4f~�fT�f��f�ʩ   uL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$�>  ���D$��~D$f��f(�f��=�  |!=2  �fT���\�f�L$�D$����f���fV��fTЗf�\$�D$���������������̃=La ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�A  ��=La t2���\$�D$%�  =�  u�<$f�$f��f���d$u�UA  ���$��  �   ��ÍT$�  R��<$t6f�<$t�-H�����=TD ��  �   ��1��  �I  �&��� u�|$ u����-��   �t���뻸   �=TD ��  �   ��1�  Z������̃=La ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�yC  ��=La t2���\$�D$%�  =�  u�<$f�$f��f���d$u�%C  ���$��  �   ��ÍT$�}  R��<$tL�D$f�<$t�-H��  �t^�   �uA������=TD ��  ��1�   �  �   �u�ԩ�� u�|$ u%   �t����-��   �"��  ���� uŃ|$ u����-���   �=TD �0  ��1�   �9  ZË�U��QSV�5 �W�5hb���5db�؉]��֋�;���   ��+��G��ruS�wF  �؍GY;�sH�   ;�s���;�rP�u��4  YY��u�C;�r>P�u��  YY��t/��P�4����hb�u�=��׉��V�ףdb�E�3�_^[�Ë�Vjj �  YY��V���hb�db��ujX^Ã& 3�^�jh`"�'  �1  �e� �u�����Y�E��E������	   �E��'  ��  Ë�U���u���������YH]�;�1u���jF  �������U��WV�u�M�}�����;�v;���  ���   r�=tb tWV����;�^_u�  ��   u������r)��$�p��Ǻ   ��r����$����$�����$��������#ъ��F�G�F���G������r���$�p��I #ъ��F���G������r���$�p��#ъ���������r���$�p��I g�T�L�D�<�4�,�$��D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�p������������E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�������$����I �Ǻ   ��r��+��$���$��� �D�l��F#шG��������r�����$���I �F#шG�F���G������r�����$����F#шG�F�G�F���G�������V�������$���I ����������������D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�����$�4�H��E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_�Ë�U��EV���F ��uc�  �F�Hl��Hh�N�;h;t� 9�Hpu�M  ��F;(8t�F� 9�Hpu��E  �F�F�@pu�Hp�F�
���@�F��^]� ��U���V�u�M��e����u�P��P  ��e�F�P�O  ��Yu��P��P  Y��xu���M����   �	��	�F�����F��u�^8M�t�E��`p��Ë�U���V�u�M�������E��u���t���   ��:�t@���u��@��t6���et��Et@���u��H�80t����   �	S�:[uH�
@B���u��}� ^t�E��`p��Ë�U����E�����Az3�@]�3�]Ë�U��QQ�} �u�ut�E�P��O  �M��E��M��H��EP�P  �E�M����Ë�U��j �u�u�u������]Ë�V����tV�Q  @PV�V�������^Ë�U��j �u�d���YY]Ë�U��j �u�����YY]Ë�U���SV�u�M�������3�;�u"�%  j^�0�}M  �}� t�E��`p���^[��9Mv�9M~�E�3���	9Ew	�~%  j"��W8Mt�U3�9M��3Ƀ:-����ˋ��6����}�?-��u�-�s�} ~�N�E�����   � � F�3�8E��E��}�u����+�]h �SV�P  ����ut�N9Et�E�G�80t/�GHy���F-��d|�jd_�� F��
|�j
_�� F�� F�LO_t�90uj�APQ�������}� t�E��`p�3������3�PPPPP��K  ̋�U���,��13ŉE��ESV�uW�}j[S�M�Q�M�Q�p�0�Q  ����u�:$  ��L  ���m�E��t���u��3Ƀ}�-��+�3Ʌ���+��M�Q�NQP3��}�-��3Ʌ�����Q��O  ����t� ��u�E�j P�u��V�u��������M�_^3�[�)����Ë�U��j �u�u�u�u�u������]Ë�U���$VW�u�M��E��  3��E�0   �Y���9}}�}�u;�u#�Z#  j^�0�K  �}� t�E�`p����  9}v؋E��� 9Ew	�$#  j"�ȋ}��E�G������  S#�3�;���   ����   �E���u�����j �u�^PSW�$�������t�}� � ��  �M�ap��  �;-u�-F�} �0����$�x�Fje��V�>  YY���U  �} ���ɀ����p��@ �;  %   �3��t�-F�]������$�x����0�F�O�����  �3���'3��u$�F0�O����� ���u�U���E��  ��F1����F�E9Uu���M܋��   �	�	��O����� �M�w;���   �U��E�   �} ~L�W#U���M�#E���� �]P  f��0����9vËM��m���E�����F�Mf�}� �E�M�}�f�}� |Q�W#U���M�#E���� �
P  f��v1�F����ft��Fu� 0H��;Et���9u��:��	�����@��} ~�uj0V�r�����u�E�8 u���} �4����$�p���W�O  3�%�  #�+E�SY�x;�r	�F+����F-������ڋ��0;�|$��  ;�rSQRP�lN  0�F�U�����;�u��|��drj jdRP�FN  0��U�F����;�u��|��
rj j
RP� N  0��U�F���]�0��F �}� t�E�`p�3�[_^�Ë�U���SVW�u���w�ٍM�N�������u#��  j^�0�G  �}� t�E��`p����   �} v׀} t;uu3��?-���f�0 �?-��u�-�s�G��V�^�J  @PVS�{����0�������} ~QV�^�pJ  @PVS�W����E����   � � ������y&�߀} u9}|�}�}������Wj0S�������}� t�E��`p�3�_^[�Ë�U���,��13ŉE��EVW�}j^V�M�Q�M�Q�p�0�4L  ����u��  �0�F  ���lS�]��u��  �0�F  ���S���;�t3Ƀ}�-����+��u�M�Q�M��QP3��}�-���P�lJ  ����t� ��u�E�j VS���N�����[�M�_3�^������Ë�U���,��13ŉE��EV�uWj_W�M�Q�M�Q�p�0�sK  ����u�  �8��E  ���   �M��t�S�]�3�K�}�-���<0���u��+ȍE�P�uQW��I  ����t� �W�E�H;������|-;E}(��t
�G��u��G��u�E�j�u���u��������u�E�jP�u���u�u������[�M�_3�^������Ë�U��E��et_��EtZ��fu�u �u�u�u�u�'�����]Ã�at��At�u �u�u�u�u�u������0�u �u�u�u�u�u�o�����u �u�u�u�u�u�o�����]Ë�U��j �u�u�u�u�u�u�Z�����]Ë�VW3��� 2���� 2����(r�_^Ë�Vh   h   3�V�kK  ����t
VVVVV��C  ^Àzuf��\���������?�f�?f��^���٭^����,��剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^����,��剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp����$����۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-���p��� ƅp���
��
�t���������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�I  ���E�f�}t�m�����������������������������������ËT$��   ��f�T$�l$é   t�   ��@��   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   �����Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t����Z��m���Z��,$Z��l������������\������   s��|���d������������T������   v��t��jh�"�x  j�J  Y�e� �u�N��t/�pD�lD�E��t9u,�H�JP�����Y�v�����Y�f �E������
   �g  Ë���j�mI  Y����̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t�����K  ��tj�K  Y�02tjh  @j��=  ��j�/  ̋�U��3��M;��t
@��r�3�]Ë��]Ë�U����  ��13ŉE�SV�uWV������3�Y�����;��l  j��O  Y���  j��O  Y��u�=hD��   ���   �6  hD�h  �xDW�@O  ������   h  ��DVSf��F�$���  ��uh�SV�O  ����t3�PPPPP�>  V��N  @Y��<v*V��N  �E4D��+�j��h�+�SP��M  ����u�h��  VW�PM  ����u������VW�<M  ����u�h  h��W�K  ���^SSSSS�y���j�� ���;�tF���tA3��G�����f9Gt@=�  r�S�����P�����P�]���@  YP�����PV���M�_^3�[�,�����j�lN  Y��tj�_N  Y��u�=hDuh�   �%���h�   ����YYË�U��E��J]�j
�(��tb3��f��QS������u����t7��$    ffAfA fA0fA@fAPfA`fAp���   HuЅ�t7����t��I f�IHu���t��3���t��IJu���t�AHu�[XË��ۃ�+�3�R�Ӄ�t�AJu���t��IKu�Z�U���W�ƃ�����   �у���te���    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tI������t��    fof�v�Ju��t$����t���v�Iu�ȃ�t	��FGIu�X^_]ú   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y����j ����,�� ��V�582�0�����u�5�J� ���V�582�4���^á42���tP�5�J� ��Ѓ42��82���tP�8��82���C  jh�"��  hx��@��u�F\��f 3�G�~�~pƆ�   CƆK  C�Fh 4j��D  Y�e� �vh�<��E������>   j�D  Y�}��E�Fl��u�h;�Fl�vl�5  Y�E������   �  �3�G�uj�C  Y�j�C  YË�VW���542��������Ћ���uNh  j��  ��YY��t:V�542�5�J� ��Ѕ�tj V�����YY���N���	V�\���Y3�W�D�_��^Ë�V��������uj�  Y��^�jh�"�  �u����   �F$��tP����Y�F,��tP����Y�F4��tP�����Y�F<��tP�����Y�F@��tP�����Y�FD��tP�����Y�FH��tP����Y�F\=�tP����Yj�@C  Y�e� �~h��tW�H���u�� 4tW�}���Y�E������W   j�C  Y�E�   �~l��t#W�4  Y;=h;t���:t�? uW�5  Y�E������   V�%���Y��  � �uj��A  YËuj��A  YË�U��=42�tK�} u'V�582�50��օ�t�542�582���ЉE^j �542�5�J� ����u�x����82���t	j P�4�]Ë�Whx��@�����u	�����3�_�V�5L�h��W��h��W��J��h��W��J��h��W��J�փ=�J �54���Jt�=�J t�=�J t��u$�0���J�8���J���5�J��J�,��82�����   �5�JP�օ���   ��  �5�J�5����5�J��J���5�J��J���5�J��J�֣�J�?  ��tc�= �h���5�J���У42���tDh  j�   ��YY��t0V�542�5�J���Ѕ�tj V����YY���N��3�@��i���3�^_Ë�U��VW3��u�v�����Y��u'9�JvV�P����  ;�Jv��������uʋ�_^]Ë�U��VW3�j �u�u�G  ������u'9�JvV�P����  ;�Jv��������uË�_^]Ë�U��VW3��u�u�G  ��YY��u,9Et'9�JvV�P����  ;�Jv��������u���_^]Ë�U��hТ�@���th��P�L���t�u��]Ë�U���u�����Y�u�T��j�?  Y�j�>  YË�V�������V��  V�3  V�����V��G  V��@  V��G  ��^Ë�U��V�u3����u���t�у�;ur�^]Ë�U��=�� th���VH  Y��t
�u���Y�G���h(�h�����YY��uTVWh���D�������Y��;�s���t�Ѓ�;�r�=pb _^thpb��G  Y��tj jj �pb3�]�j h�"�[  j�>  Y�e� 3�@9�J��   ��J�E��J�} ��   �5hb�5 ��֋؉]Ѕ�th�5db�֋��}ԉ]܉}؃��}�;�rK����9t�;�r>�7�֋��r�������5hb�֋��5db��9]�u9E�t�]܉]ЉE؋��}ԋ]���E�,��}�8�s�E� ��t�ЃE����E�<��}�@�s�E�� ��t�ЃE����E������    �} u)��J   j�<  Y�u�����} tj�<  Y��m  Ë�U��j j�u������]�jj j ������Ë�U���x����u�����Yh�   ����̋�U���LV�E�P�d�j@j ^V����YY3�;�u����  ��   �`a�5Ta;�s6���H��f�@� 
�Hf�@ 
�@!
�H3�H/�5`a��@�P���   ;�r�SWf9M��  �E�;��  ����E�þ   �E�;�|��9Ta}k�daj@j �����YY��tQ�Ta ��   �;�s1���H���` �`��`3 f�@� 
f�@ 

�@/ ���@΍P�;�r҃�9Ta|���Ta3���~r�E�� ���t\���tW�M��	��tM��uP�`���t=����������4�`a�E�� ��E�� �Fh�  �FP�\�����   �F�E�G�E�;�|�3ۋ���5`a����t���t�N��q�F���uj�X�
�C�������P� ������tB��t>W�`���t3%�   �>��u�N@�	��u�Nh�  �FP�\���t,�F�
�N@�����C���h����5Ta�X�3�_[^�Ã������VW�`a���t6��   ;�s!�p�~� tV�h����@   �N�;�r��7������' Y����`b|�_^Ã=lb u�a+  V�5\DW3���u����   <=tGV�M3  Y�t���u�jGW�������YY�=�J��tˋ5\DS�3V�3  �>=Y�Xt"jS����YY���t?VSP�3  ����uG���> u��5\D�A����%\D �' �`b   3�Y[_^��5�J�����%�J �����3�PPPPP�#/  ̋�U��Q�MS3�V���U�   9Et	�]�E��E��>"u3�9E��"��F�E��<���t��B�U���PF�C  Y��t��} t
�M��E�F�U�M��t2�}� u��� t��	u���t�B� �e� �> ��   �< t<	uF��N��> ��   �} t	�E�E��3�C3��FA�>\t��>"u&��u�}� t�F�8"u���3�3�9E����E����tI��t�\B���u�U���tU�}� u< tK<	tG��t=��P��t#�B  Y��t��M�E�F��M��E���B  Y��tF���UF�V�����t� B�U��M�����E^[��t�  ��Ë�U���S3�VW9lbu��(  h  ��JVS��K�l��xb�5�J;�t�E�8u�u��U��E�PSS�}��
����E���=���?sJ�M���sB�����;�r6P�������Y;�t)�U��E�P�WV�}�������E���H��J�5�J3�����_^[�Ë�U���SV�x���3�;�u3��wf93t��f90u���f90u�W�=t�VVV+�V��@PSVV�E��׉E�;�t8P�;���Y�E�;�t*VV�u�P�u�SVV�ׅ�u�u��4���Y�u�S�p��E��	S�p�3�_^[�Ë�V�"�"W��;�s���t�Ѓ�;�r�_^Ë�V�"�"W��;�s���t�Ѓ�;�r�_^�j h   j �|�3Ʌ�����K����5�K����%�K �������h��d�5    �D$�l$�l$+�SVW��11E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q�������̋�U���S�]V�s35�1W��E� �E�   �{���t�N�38�����N�F�38�����E�@f�  �M�U�S��[�E�M���t_�I �[�L��D��E�� �E���t���t6  �E���x@G�E��؃��u΀}� t$����t�N�38�����N�V�3:�~����E�_^[��]��E�    �ɋM�9csm�u)�=Pa t hPa�>  ����t�UjR�Pa���M�U�6  �E9Xth�1W�Ӌ��6  �E�M��H����t�N�38������N�V�3:������E��H���5  �����9S�O���h�1W����5  ������U��V����������2  �N\�U��W9t�����   ;�r���   ;�s9t3���t�P��u3���   ��u�` 3�@��   ����   �MS�^`�N`�H����   j$Y�~\�d9 �����   |� �~d=�  �u	�Fd�   �~=�  �u	�Fd�   �n=�  �u	�Fd�   �^=�  �u	�Fd�   �N=�  �u	�Fd�   �>=�  �u	�Fd�   �.=�  �u	�Fd�   �=� �u	�Fd�   �=� �u�Fd�   �vdj��Y�~d��` Q��Y�^`[���_^]Ë�U��csm�9Eu�uP����YY]�3�]Ë�U�����1�e� �e� SW�N�@��  ��;�t��t	�У�1�eV�E�P����u�3u����3���3����3��E�P����E�3E�3�;�u�O�@����u��G  ����5�1�։5�1^_[�Ë�U��E3�;̀2tA��-r�H��wjX]Ë̈́2]�D���jY;��#���]�������u��3Ã���~�����u��3Ã�Ë�U��V������MQ�����Y�������0^]Ë�U��E��K]Ë�U���5�K� ���t�u��Y��t3�@]�3�]�j
�(��La3������������U�������$�~$�   ��fD$f%0�f@�fW�f8���fs�,f~����    f������� #�- � =�  ��   �YɁ���  �\��Q�fT׃���� �  fU��fV�f($������X��\��Y��Y��Y����X��^�f=�f-غ�\�fs�?��fs�?�Y�fp�Df5��Y��Y���fW��Y��Y��X��Y��X�fp���X��X��X�fD$�D$���-�  ��C�  �Y��\��Q�f��fs�fT=кfs���f%@����\��Y��X��\��Y���fT�fs�f��fVՁ���  ��Y<����Y�f(���Y��Y��\��X��\��X�f-غ�\��X�f��^�f�f\ՠ����Y�%�   ���Y��Y΃��Y��Y��X�f���Y��X�f���X�fp���\��X�fV�fD$�D$����;  = 8  sjf�f(5�f�f( �f(%�fY���fY�fY�fY����Y�fX�fY��Y�fX�fY�fp���X��X�fD$�D$���-�;  ���O  �Y��\��Q�f��fT=��fp�DfT����f%@����\��Y��X��Y��\����Y��Y��\��\��X��\�f(�fp���\��X�fp���X��Y��X�fp���^�f( �f(- �f(�fY���fY�fY�% �  �Y�fY�fX�f(��Y�fY�f(���Y�fX�fp���Y��fY��X�fW�fp���Y�fp���X���f���\��X��X��X��\��\��\��\�fV�fD$�D$����� = � ��   f~�fs� f~�����  �?+���� ��   fT$f~�fs� f~с��������  ��� ��   fW�fW���  f���Y��=   ��fD$�T$�ԃ��T$���T$�$�	  fD$����fD$�D$���f0�f��f���X�fU�fV���fD$�D$���fD$fW��Xƺ�  �t���fD$fW�����f�����  �����  r�X�fV��Y�fD$�D$���U�������$�~$�   ��fD$f%@�fP�fW�fH���fs�,f~����    f������� #�- � =�  ��   �YɁ���  �\��Q�fT׃���� �  fU��fV�f($������X��\��Y��Y��Y����X��^�f��f-���\�fs�?��fs�?�Y�fp�Df5���Y��Y���fW��Y�f\%���Y��X��Y��\�fp���X��\��\�fD$�D$���-�  ��A�-  fs�&fs�&f��fU��\����Y��X�fV��\��Y����\��Q�%�   ������fT�fs�f��fV�fn�fp� ����  ��Y<����Y��Y��Y��\�fT���X��\��X�f-���\��X�f���^�f��fXՀ����Y��Y��Y΃��Y��Y��X�f���Y��X��X�% �  f����fp���X��\��X��X��X�fW�fD$�D$����;  = 8  ��   f�f(5 �f�f(�f(% �fY�f(-����fY�fY�fY����Y�fX�fY��Y�fX�fp��fY�fp���\�fp���\��\��\��\��\��X�fD$�D$���-�;  ����   fW�fT=@�f%X�f( ��Y�f(��\�f( �fp�D�Q�fY�fp�Df��fY�fX�f��fY�����Y�fX�fp�D�Y�fT��fY�fT�fp�D�\��X��Y��\��\��Y�fp���\��^��fX�fY�fp���X�% �  f��fp���X��X��X��X�fW�fD$�D$����� = � ��   f~�fs� f~�������  �?+���� ��   fT$f~�fs� f~с��������  ��� ��   fW�fW���  f���Y��:   ��fD$�T$�ԃ��T$���T$�$�  fD$����fD$�D$���f������fn�fp� f��f��fT�fT��X�fD$�D$���f��f���X�fD$�D$���fW��Xƺ�  �J���������������U�������$�~$�   ��fD$f��f%�f-00f=��B  f���Y�f���-��X�f���\�f(���Y�fɁ�v ����?f(-��������fY��\��Y���\�fxf����\�fY�f\�f(5���Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-���Y fX5��fY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X΃��X�fd$�D$���+f��f%�f����f ��\�fL$�D$��������I ����U�������$�~$�   ��fD$f��f%�f-00f=��B  f���Y�f���-��X�f���\�f(���Y�fɁ� v ����?f(-p��@����fY��\��Y���\�fxf����\�fY�f\�f(5P��Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-`��Y fX5@�fY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X΃��X�fd$�D$���I��f��f=�u�Y��fD$�D$���f���Y��\��Y��fD$�D$����������U���(3��E��E�9Lt�5Ha� ����&�M��   V;���  ��  ���  �  jZ+���   I��   ����   I��   ����   ItN��	�  �E�   �Eܜ��M��M�u�]���M��]�Q��]���Y����  �L���� "   ��  �Eܘ��M��M�u�]���M��]�Q��E�   �]���Y�  �E�   �Eܘ���Eܐ��M�u��M�]���]���?  �U��Eܐ��W����E܌��ΉU��E܌��?����Eܜ��q�����tWItHIt9It ��t���  �E܄���E�|���Eܜ��M��u��u����Eܜ��c����E�   �������E���   �E�   �E�t��������������   �$� ��E܌���Eܐ���Eܘ���E�l���E�d��t����E�\��h����E�T��\����E�P���E�L���E�H��M��u�M����M�]���]�M��]�Q�E�   ��Y��u����� !   �E��^�Ð\�e�n�w��������������������U��QQSV���  V�5�3�3  �EYY�M�ظ�  #�QQ�$f;�uU�1  YY��~-��~��u#�ESQQ�$j�/0  ���tVS��2  �EYY�f�ES�ؑ���\$�E�$jj�A�1  �]��E�Y�EY������DzVS�2  �E�YY�"�� u��E�S���\$�E�$jj�0  ��^[������U�������$�~<$�   ���~|$f�f(�fT��f/����  �U  f/��snf/����  f(�fY�f(�fY�f(-��fY�fX-p�fY�fX-`�fY�fX-P��Y�f(�f���X��Y��\�f�|$�D$�f/����   f(�fY�f(�fY�f(-@�fY�fX-0�fY�fX- �fY�fX-�fY�fX- �fY�fX-��fY�fX-��fY�fX-���Y�f(�f���X��Y��\�f�|$�D$��~�fW�f/��sO�~���~-���~��X�fs�,f��f~؍@�~,����~��\��Y��X���^�f���   �~��~���^�f��~����~$���f(�fY�f(�fY�f(-��fY�fX-p�fY�fX-`�fY�fX-P��Y�f(�f���X��Y��\��\��\�fV�f�D$�D$�f/��u�D$�f/��s���������$�$���D$��������D$��~��~��fT�f.�z�D$���������ú�  ���T$�ԃ��T$�T$�$�u������D$Ð����U�������$�~$�   ��fD$�    f(�f�fs�4f�� f(��f(P�f(% �f(5�fT�fV�fX�f�� %�  f(���f(���fT�f\�fY�f\��X�fY�f(�fXƁ��  �����  ��   ���  ��*�f���
��   �    �� D�f(��f(�f(��fY�fY�fX�f(���Y�f(- �fY�f(�0�fT�fX�fX�fY��Y�fX�f(�f�fY˃�f(�f��X��X��X�fD$�D$���fD$f(`���� f�� �� wH���t^���  wlfD$f(��f(P�fT�fV���� f�� �� t���ú�  �OfP��^�f���   �4fp��Y�������/��������  ���  s:fW��^ɺ   ��fL$�T$�ԃ��T$���T$�$�1����D$���fT$fD$f~�fs� f~с��� ��� t���  릍d$ ƅp����
�u;�����ƅp����2������+  ������a���t������@u��
�t���B����F  �t2��t��������8�������������-��ƅp����������ݽ`������a���Au����ƅp������-���
�uS��������
�u�����������   ����
�u���u
�t���ƅp����-����u�
�t��������������8���X��ݽ`������a���u���-��
�t���ƅp����g��������-��ƅp����
�u����-��������-��ٛݽ`������a���Au�������ݽ`������a���������ݽ`�������������ٛ���u���"������ٛ���t�   ø    ���   ��V��t��V���$���$��v�v,  ���f���t^��t�S���Ë�U��} u������    ��  ���]��uj �5�K���]Ë�U��� �e� Wj3�Y�}��9Eu�����    �~  ����x�MV�u��t��u�����    �Z  ����S�����E�;�w�M��u�E��u�E�B   �u�u�P�u���.  ������t�M�x�E��  ��E�Pj �,  YY��^_�Ë�U���uj �u�u�u�<�����]Ë�U���(  �M�M�M�M�5 M�=�Lf�(Mf�Mf��Lf��Lf�%�Lf�-�L�� M�E �M�E�M�E�$M�������`L  �M�L�L	 ��L   ��1��������1����������XLj��9  Yj ���hL�����=XL uj�9  Yh	 ����P������������U��W�}3�������ك��E���8t3�����_��-�  t"��t��tHt3�ø  ø  ø  ø  Ë�VW��h  3��FWP�����3��ȋ��~�~�~����~���� 4���F+ο  ��@Ou���  �   ��@Nu�_^Ë�U���  ��13ŉE�SW������P�v����   ����   3�������@;�r�����ƅ���� ��t0���������;�w+�@P������j R�:������C����u�j �v�������vPW������Pjj �<;  3�S�v������WPW������PW�vS��9  ��DS�v������WPW������Ph   �vS��9  ��$3���E������t�L���������t�L ��������  ���  @;�r��R��  ǅ��������3�)�������������  ЍZ ��w
�L�Q ���w�L �Q����  A;�rƋM�_3�[�,�����jh#�t���������� 9�Gpt�l t�wh��uj �M���Y�������j�o  Y�e� �wh�u�;5(8t6��tV�H���u�� 4tV衫��Y�(8�Gh�5(8�u�V�<��E������   뎋u�j�5  YË�U���S3�S�M������,O���u�,O   ���8]�tE�M��ap��<���u�,O   ����ۃ��u�E��@�,O   ��8]�t�E��`p���[�Ë�U��� ��13ŉE�S�]V�uW�d�����3��};�u������3��  �u�3�9�08��   �E��0=�   r����  �t  ����  �h  ��P������V  �E�PW������7  h  �CVP�]���3�B���{�s9U���   �}� ��   �u�����   �F����   h  �CVP�����M��k�0�u���@8�u��+�F��t)�>����E���,8D;�FG;�v�}���> uЋu��E����}��u�r�ǉ{�C   �i���j�C�C��48Zf�1f�0����Ju������������L@;�v����~� �0����C��   �@Iu��C�����C�S��s3��ȋ�����{����95,O�T�������M�_^3�[�#�����jh0#�k����M���������}�������_h�u�q����E;C�W  h   ����Y�؅��F  ��   �wh���# S�u����YY�E�����   �u��vh�H���u�Fh= 4tP�y���Y�^hS�=<����Fp��   � 9��   j��  Y�e� �C�<O�C�@O�C�DO3��E��}f�LCf�E0O@��3��E�=  }�L�� 6@��3��E�=   }��  ��(7@���5(8�H���u�(8= 4tP�����Y�(8S���E������   �0j�f  Y��%���u �� 4tS芧��Y�(����    ��e� �E��#���Ã=lb uj��V���Y�lb   3�Ë�U��SV�5<�W�}W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{�$9t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��_^[]Ë�U��W�}����   SV�5H�W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{�$9t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��^[��_]Ë�U��SV�u���   3�W;�to=�=th���   ;�t^9uZ���   ;�t9uP�������   �;8  YY���   ;�t9uP�ȥ�����   �7  YY���   谥�����   襥��YY���   ;�tD9u@���   -�   P脥�����   ��   +�P�q������   +�P�c������   �X��������   =(9t9��   uP�3  ���   �/���YY�~P�E   ��$9t�;�t9uP�
���Y9_�t�G;�t9uP����Y���Mu�V����Y_^[]Ë�U��W�}��t;�E��t4V�0;�t(W�8�j���Y��tV������> Yu���:tV�s���Y��^�3�_]�jhP#������3����� 9�Fpt"�~l t�����pl��uj �����Y�������j��  Y�e� �5h;��lV�Y���YY�E��E������   �j��
  Y�u�Ë�U��E�HO]Ë�U���(  ��13ŉE�S�]W���tS�/  Y������ jL������j P�ڜ����������������0�����������������������������������������������f������f������f������f������f������f��������������E�M������ǅ0���  �������I��������M�������M���������������j �����������P�����u��u���tS�.  Y�M�_3�[������Ë�Vj� �Vj�������V���P���^Ë�U���5HO� ���t]���u�u�u�u�u�����3�PPPPP�������Ë�U����u�M�������E����   ~�E�Pj�u�5  ������   �M�H���}� t�M��ap��Ë�U��=Q u�E�X;�A��]�j �u����YY]Ë�U���SV�u�M��y����]�   ;�sT�M胹�   ~�E�PjS�!5  �M������   �X����t���   ��   �}� t�E��`p����   �E胸�   ~1�]�}�E�P�E%�   P�x5  YY��t�Ej�E��]��E� Y������� *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QV�p�E�P�(.  ��$���o������E�t	�M�����}� t�M��ap�^[�Ë�U��=Q u�E�H���w�� ]�j �u�����YY]Ë�U���(��13ŉE�SV�uW�u�}�M��'����E�P3�SSSSW�E�P�E�P�?  �E�E�VP��4  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�0����Ë�U���(��13ŉE�SV�uW�u�}�M������E�P3�SSSSW�E�P�E�P��>  �E�E�VP�z9  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[舩���������������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+�Ë�U��UVW��t�}��u�a���j^�0�%������3�E��u����+���@��tOu��u� �+���j"Y�����3�_^]Ë�U��MS�YV�u3�;�u����j^�0��������   9Ev�U�;�~��@9Ew�����j"Y�����W�~�0�ǅ�~���t��C�j0Y�@J���M�  ��x�;5|�� 0H�89t�� �>1u�A�W�v���@PWV�]�����3�_^[]Ë�U��Q�M�AS����% �  V��  #�W�E�A�	���   �%�� �u���t;�t�� <  �(��  �$3�;�u;�u�Ef�M�P��B��<  �U����������U��E����������Ɂ���  ��P��t�M�_^f�H[�Ë�U���0��13ŉE��ES�]V�E�W�EP�E�P�"���YY�E�Pj j���uЋ���f��B  �u܉C�E��E��C�E�P�uV�������$��u�M�_�s^��3�[諦����3�PPPPP�������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��j�����YË�U��E�M%����#�V�u������t$��tj j �QK  YY������j^�0�������P�u��t	�-K  ���$K  YY3�^]Ë�S��QQ�����U�k�l$���   ��13ŉE��C�V�s�HW��x���tRHtCHt4Ht%HtFHHtH��   ǅ|���   �9�   �   ǅ|���   �"ǅ|���   �ǅ|���   �
ǅ|���   Q�~W��|����y  ����uI�C��t��t��t�e����M��F����]����M�W�NQP��|�����x���P�E�P�	  ��h��  ��x����  �>YYt�=�< uV�  Y��u�6��  Y�M�_3�^�������]��[Ë�VW3��PO�<�t;u��p;�8h�  �0���\���tF��$|�3�@_^Ã$�p; 3����S�h�V�p;W�>��t�~tW��W�m����& Y�����<|ܾp;_���t	�~uP�Ӄ����<|�^[Ë�U��E�4�p;���]�jhp#����3�G�}�3�9�Ku����j�;���h�   �����YY�u�4�p;9t���mj輿��Y��;�u�o����    3��Pj
�X   Y�]�9u+h�  W�\���uW蜘��Y�:����    �]���>�W聘��Y�E������	   �E������j
�)���YË�U��EV�4�p;�> uP�#���Y��uj����Y�6���^]��������������SVW�T$�D$�L$URPQQh@d�5    ��13ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�L  �   �C�L  �d�    ��_^[ËL$�A   �   t3�D$�H3�芡��U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j��K  3�3�3�3�3���U��SVWj Rh�Q�,f  _^[]�U�l$RQ�t$������]� ��U��E��P��P��P��P]Ë�U��E���V9Pt��k�u��;�r�k�M^;�s9Pt3�]��5�P� ��j h�#�����3��}�}؋]��Kt��jY+�t"+�t+�tY+�uC�p������}؅�u����T  ��P��P�U�w\���]���Y�p��Q�Ã�t2��t!Ht�����    �Z���빾�P��P���P��P�
��P��P�E�   P� ��E�3��}���   9E�uj����9E�tP�.���Y3��E���t
��t��u�O`�MԉG`��u>�Od�M��Gd�   ��u,�x��M܋|�x�9M�}�M�k��W\�D�E����-�����E������   ��u�wdS�U�Y��]�}؃}� tj ����Y�S�U�Y��t
��t��u�EԉG`��u�EЉGd3�����Ë�U���$��13ŉE��ES�E��EVW�E�訶���e� �=�P �E�u}h0��Ȑ�؅��  �=L�h$�S�ׅ���   �5�P��h�S��P��P��h �S��P��P��h��S��P��P�֣ Q��th��S��P�֣�P��P�M�5 �;�tG9 Qt?P���5 Q���֋؅�t,��t(�ׅ�t�M�Qj�M�QjP�Ӆ�t�E�u	�M    �3��P;E�t)P�օ�t"�ЉE��t��P;E�tP�օ�t�u��ЉE��5�P�օ�t�u�u��u��u����3��M�_^3�[�y����Ë�U��V�uW��t�}��u�����j^�0������_^]ËM��u3�f��݋�f�: t��Ou��t�+��f�
��f��tOu�3���u�f�����j"Y���몋�U��US�]VW��u��u9Uu3�_^[]Å�t�}��u�\���j^�0� ������݅�u3�f��ЋM��u3�f��ԋ��u��+��f���f��t'Ou��"��+��f���f��tOtKu��u3�f����y���3����u�MjPf�DJ�X�d���f������j"Y����j�����U��Ef���f��u�+E��H]Ë�U��V�uW��t�}��u����j^�0�P�����_^]ËE��uf��ߋ�+��f���f��tOu�3���u�f��L���j"Y���뼋�U��M��x��~��u�dD]ádD�dD]������    ��������]Ë�U��E��t���8��  uP�C���Y]Ë�U��M��tj�3�X��;Es������    3�]��MV���uF3����wVj�5�K����u2�= L tV�����Y��uҋE��t�    3���M��t�   ^]Ë�U��} u�u����Y]�V�u��u�u蘐��Y3��MW�0��uFV�uj �5�K�̐����u^9 Lt@V�a���Y��t���v�V�Q���Y������    3�_^]����������P����Y������������P�z���Y�����jh�#�s���賳���@x��t�e� ���3�@Ëe��E������ĭ�������h�$���QË�U��E�Q]������̋�U��M�MZ  f9t3�]ËA<��8PE  u�3ҹ  f9H��]�����������̋�U��E�H<��ASV�q3�W�D��t�}�H;�r	�X�;�r
B��(;�r�3�_^[]������������̋�U��j�h�#h��d�    P��SVW��11E�3�P�E�d�    �e��E�    h   �*�������tT�E-   Ph   �P�������t:�@$���Ѓ��E������M�d�    Y_^[��]ËE�3ҁ9  ���Ëe��E�����3��M�d�    Y_^[��]Ë�U����u�M������E�M�U�Tu�} t�M����   �A#E�3���t3�@�}� t�M��ap��Ë�U��jj �uj ������]�3�Ë�U��E�MSVW3��x�E3ۉx�EC�x��t�E	X�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ��u��E����3H��1H��E���3H��1H��E����3H��1H��E����3H��1H��E����3H#�1H�  ��t�M�I�t�M�I�t�M�I�t�M�I� t�E	X��   #�t5=   t"=   t;�u)�E��!�E���������E��������E� ���   #�t =   t;�u"�E� ���E�������E�������E�M��3���� 1�E	X 9} �E�}t&�` �E� �E�X�E	X`�E�``���E�XP�4�H �����H �E� �E�X�E	X`�E�H`�����H`��E�XP�c  �EPSj �u�А�M�At�&��At�&��At�&��At�&�Yt�&ߋ��3�+ú����t/HtHtHu(�   � �%����   ���%����   ��!�����+�tHtHu!��#�   �	�#�   �9] t�AP���AP�_^[]Ë�U��j �u�u�u�u�u�u������]Ë�U����ESV3ۋ���C�u��t�]tS�  Y����  �t�Etj�y  Y����x  ����   �E��   j�W  �EY�   #�tT=   t7=   t;�ub��M�����=��{L�H��M�����{,��=�2��M�����z��=���M�����z��=���=��������   ���   �E��   3��t��W�}���������D��   ��E�PQQ�$�  �M��]�� �����������}�E������S���]�����Au���3ҋE����f�E����;�}"+��]�t��u���m�]�t�M�   ��m�Hu���t�E����]��E�����_��tj�   Y�e���u��Et�E tj ��  Y���3���^��[�Ë�U��}t~�}衾��� "   ]�蔾��� !   ]Ë�U��E� tj��t3�@]ètj��tjX]������]Ë�U��� 3��Ř<;Mtd@��|�3��E��t^�E�E�E�E�E�E��EV�u�E�E �E��E$h��  �u(�u��E���  �E�P�S�������uV�,���Y�E�^�ËŜ<�h��  �u(�  �u�����E ���Ë�U��=�< u(�u�E���\$���\$�E�$�uj�/�����$]��}���h��  �u� !   �\  �EYY]Ë�S��QQ�����U�k�l$���   ��13ŉE��s �CP�s��������u#�e��P�CP�CP�s�C �sP�E�P�j������s�o������=�< u+��t'�s �C���\$���\$�C�$�sP�q�����$�P�����$��  �s �  �CYY�M�3�������]��[Ë�U��QQ�E���]��E��Ë�U��QQ�E�E�M�]��  �����  �f�E��E��Ë�U��3ҁ}  �u
9Uu3�@]Á}  ��u
9UujX]�f�M��  V��f#�^f;�uj���  f;�u�E�� u9Utj��3�]Ë�U���E������������Dz3��   �E3ɩ�  uk�E�� u9Mt]�]��������Au3�@�3���e�E   �t�M�eJ�Et�V���  f!u^;�t	� �  f	E�EQQQ�$��������&Q���EQQ�$������U�����  �����  �E�]Ë�U��Q��}��E��Ë�U��Q�}����E��Ë�U��Q��}��E�M#M��f#E�f����E�m�E��Ë�U��QQ�M��t
�-�=�]���t����-�=�]�������t
�-�=�]����t	�������؛�� t���]����jh�#�I���3�9tbtV�E@tH9�=t@�E��U�.�E� � =  �t
=  �t3��3�@Ëe�%�= �e��U�E�������e��U�)���Ë�U��QQ�EQQ�$�9  YY��uL�EQQ�$�Y����EY��Y����Dz1�EQ�8�Q�]��E��$�2����E�Y��Y����DzjX��3�@��3��Ë�U���EV�  ���3�3��  ��9Eu:9Uuz��������z������=��   ��������A�E��   ������   9Mu@9Uu;��������z�������   ������A�Eu��=�   ��=3�F�   ��9Eu(9Uu}���U�����w����U����A�Et^�����X9MuU9UuP�EQQ�$������Y�UY������z����=��u!����U����Au��u����=�����E���^]Ë�U��QV�uV�+D  �E�FY��u�d���� 	   �N ����/  �@t�I���� "   ��S3ۨt�^���   �N�����F�F�����F�^�]��  u,�B  �� ;�t��A  ��@;�u�u�A  Y��uV�CA  Y�F  W��   �F�>�H��N+�I�N;�~WP�u�?@  ���E��M�� �F����y�M���t���t�����������`a��@2�@ tjSSQ�8  #����t%�F�M��3�GW�EP�u��?  ���E�9}�t	�N �����E%�   _[^���A@t�y t$�Ix��������QP�v���YY���u	��Ë�U��Q�C@V����E�t�{ u�E�>�' �} ~0�E� �M�������E�>�u�?*u�˰?�~����} Ճ? u�E��^�Ë�U���  ��13ŉE�S�]V�u3�W�}�u����������������������������������������������������������������������������u+�����    ����������� t
�������`p�����7  �F@u^V�A  Y�@2���t���t�ȃ��������`a����A$u����t���t�ȃ������`a����@$��q���3�;��g��������������������������������
  C3�������9������y
  �B�<Xw��������3�����j��Y������;�� 
  �$��?���������������������������������������������	  �� tJ��t6��t%HHt����	  �������	  �������	  �������	  �������   �	  �������	  ��*u,����������������;��l	  �������������Z	  ������k�
�ʍDЉ������?	  �������4	  ��*u&����������������;��	  ��������		  ������k�
�ʍDЉ�������  ��ItU��htD��lt��w��  ������   ��  �;luC������   �������  �������  ������ �  �<6u�{4u�������� �  �������p  <3u�{2u������������������N  <d�F  <i�>  <o�6  <u�.  <x�&  <X�  ������!�����������P��P�b  Y��������Yt"�����������������C������������������������������  ��d��  �X  ��S��   tL��AtHHt$HHtHH��  �� ǅ����   �������V  ������0  ��   ������   �   ������0  u
������   ���������u������������  ����������������  ��u��=������������ǅ����   ��  ��X�"  HHt+���  HH��  ��������������  ������t0�G�Ph   ������P������P��>  ����tǅ����   ��G�������ǅ����   �������������|  �����������t;�H��t4������   � ������t�+���ǅ����   �7  !������,  ��=������P�����Y�  ��p�=  �%  ��e�  ��g��   ��it|��nt.��o��  �������������ǅ����   tl������   �`�������������p��\<  ���b��������� tf������f���������ǅ����   �>  ������������@ǅ����
   �������� �  ��  ��W���  ������������@�������   ������������9�����}ǅ����   �ju��gucǅ����   �W9�����~�������������   ~=��������]  V�ߠ��������Y��������t���������������
ǅ�����   ��5 ����������G�������������P��������������������P������������SP�52���Ћ���������   t������ u������PS�5$2����YY������gu��u������PS�5 2����YY�;-u������   C������S�����ǅ����   �������*��s�n���HH�X�������  ������ǅ����'   �������ǅ����   �2���������Qƅ����0������ǅ����   ������   �������� t��������@t�G���G����G���@t��3҉�������@t��|��s����ځ�����   ������ �  ����u3�9�����}ǅ����   ���������   9�����~���������u!������u����������������t-�������RPWS��*  ��0�������؋���9~������N뽍E�+�F������   ������������tb��t�΀90tW�������������0@�?If90t����u�+��������(��u��=�������������I�8 t@��u�+����������������� ��  ��������@t5��   t	ƅ����-���t	ƅ����+���tƅ���� ǅ����   ������+�����+�������������u%���������������� O�0����������t���������������������������P�������2���������YYt.������u%��������������˰0O������������t��ヽ���� ������tu��~q�������������������Pj�E�P������P����8  ����u69�����t.�������������������E�P���������������� YYu��#��������������P�������������]���YY������ |2������t)�������������������� O������������t��߃����� t�������Uu�������� Y���������������t���������������r��������� t
�������`p��������M�_^3�[����Ðm7l5�5�5F6Q6�6�7�%Da Ë�U�����13ŉE��US3�VW;�~�E��I8t@;�u������+�H;�}@�E�]�9]$u�E� �@�E$�5ؐ3�9](SS�u���u��   P�u$�֋��}�;�u3��R  ~Cj�3�X����r7�D?=   w�4)  ��;�t� ��  �P�s��Y;�t	� ��  ���E���]�9]�t�W�u��u�uj�u$�օ���   �5ԐSSW�u��u�u�։E�;���   �   �Mt)�E ;���   9E���   P�uW�u��u�u���   �}�;�~Bj�3�X����r6�D?;�w�z(  ��;�th���  ���P��r��Y;�t	� ��  �����3�;�t?�u�W�u��u��u�u�օ�t"SS9] uSS��u �u�u�WS�u$�t��E�W����Y�u������E�Y�e�_^[�M�3��
}���Ë�U����u�M��l����u(�E��u$�u �u�u�u�u�uP�������$�}� t�M��ap��Ë�U��QQ��13ŉE�S3�VW�]�9]u�E� �@�E�5ؐ3�9] SS�u���u��   P�u�֋�;�u3��~<�����w4�D?=   w�8'  ��;�t� ��  �P�q��Y;�t	� ��  ���؅�t��?Pj S�k����WS�u�uj�u�օ�t�uPS�u�ܐ�E�S�y����E�Y�e�_^[�M�3���{���Ë�U����u�M��?���u$�E��u�u�u�u�uP��������}� t�M��ap��Ë�U��V�u���c  �v�jq���v�bq���v�Zq���v�Rq���v�Jq���v�Bq���6�;q���v �3q���v$�+q���v(�#q���v,�q���v0�q���v4�q���v�q���v8��p���v<��p����@�v@��p���vD��p���vH��p���vL��p���vP��p���vT��p���vX�p���v\�p���v`�p���vd�p���vh�p���vl�p���vp�p���vt�p���vx�xp���v|�pp����@���   �bp�����   �Wp�����   �Lp�����   �Ap�����   �6p�����   �+p�����   � p�����   �p�����   �
p�����   ��o�����   ��o�����   ��o�����   ��o�����   ��o�����   ��o�����   �o����@���   �o�����   �o�����   �o�����   �o�����   �o�����   �xo�����   �mo�����   �bo�����   �Wo�����   �Lo�����   �Ao�����   �6o�����   �+o����   � o����  �o����  �
o����@��  ��n����  ��n����  ��n����  ��n����  ��n����   ��n����$  �n����(  �n����,  �n����0  �n����4  �n����8  �n����<  �xn����@  �mn����D  �bn����H  �Wn����@��L  �In����P  �>n����T  �3n����X  �(n����\  �n����`  �n����^]Ë�U��V�u��tY�;�=tP��m��Y�F;�=tP��m��Y�F;�=tP��m��Y�F0;>tP�m��Y�v4;5>tV�m��Y^]Ë�U��V�u����   �F;�=tP�m��Y�F;�=tP�om��Y�F;�=tP�]m��Y�F;�=tP�Km��Y�F;�=tP�9m��Y�F ;�=tP�'m��Y�F$;�=tP�m��Y�F8;>tP�m��Y�F<;>tP��l��Y�F@;>tP��l��Y�FD;>tP��l��Y�FH; >tP�l��Y�vL;5$>tV�l��Y^]Ë�U���S�u�M�� z���]�C=   w�E苀�   �X�u�]�}�E�P�E%�   P�o   YY��t�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�p�E�PQ�E�P�E�jP�X����� ��u8E�t�E��`p�3���E�#E�}� t�M��ap�[�Ë�U����u�M��iy���E�M����   �A% �  �}� t�M��ap��Ë�U��j �u����YY]Ë�U���8��13ŉE��E�M�M��H
S�ف� �  �MȋH�M��H� ���  ���?  ��W�M�E������u'3�3�9\��u@��|�3��  3��}�j�X�  �e� V�u��}䥥��=@>O�G�������W��  ��]ԉE�yJ���B�t��j3�Y+�@���MЅ��   �E؃�����҅T����|�� u@��|��n�ǙjY#������  �yO���G�e� +�3�B��L���9��}��99}�r"9U����t+�e� �L����z�}�;�r��s�E�   H�U���M�yщM܋MЃ����jY!�E�@;�}
�|��+�3��}� tC�<>��+@>;�}3��}𫫫�	  ;��  +Eԍu�ȍ}𥙃�¥������  ��yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�5@>N�F�������V��  ��E�yJ���BjY+�3�B��\���Mԅ��   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e� 3�+�B��L���1�<;�r;�s�E�   �9�M����t�L����r3�;�r��s3�G�1��HyދMԃ����!�E�@��}jY�|��+�3��D>�A���Q����  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�j3�X�S  �D>;8>��   3��}𫫫�M�   �����������  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�L>8>3�@�   L>�e��������������  �yJ���B�e� �e� ��������E�    )U��֋M��|����#ΉMԋ���M�}؉|���}ԋM����E��}��}�|Ћ�j���M�Z+�;�|�1�t����d�� ��Jy�3�^jY+D>��M���Ɂ�   �ًH>]���@u�M̋U�Y��
�� u�M̉�M�_3�[�kp���Ë�U���8��13ŉE��E�M�M��H
S�ف� �  �MȋH�M��H� ���  ���?  ��W�M�E������u'3�3�9\��u@��|�3��  3��}�j�X�  �e� V�u��}䥥��=X>O�G�������W��  ��]ԉE�yJ���B�t��j3�Y+�@���MЅ��   �E؃�����҅T����|�� u@��|��n�ǙjY#������  �yO���G�e� +�3�B��L���9��}��99}�r"9U����t+�e� �L����z�}�;�r��s�E�   H�U���M�yщM܋MЃ����jY!�E�@;�}
�|��+�3��}� tC�T>��+X>;�}3��}𫫫�	  ;��  +Eԍu�ȍ}𥙃�¥������  ��yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�5X>N�F�������V��  ��E�yJ���BjY+�3�B��\���Mԅ��   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e� 3�+�B��L���1�<;�r;�s�E�   �9�M����t�L����r3�;�r��s3�G�1��HyދMԃ����!�E�@��}jY�|��+�3��\>�A���Q����  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�j3�X�S  �\>;P>��   3��}𫫫�M�   �����������  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�d>P>3�@�   d>�e��������������  �yJ���B�e� �e� ��������E�    )U��֋M��|����#ΉMԋ���M�}؉|���}ԋM����E��}��}�|Ћ�j���M�Z+�;�|�1�t����d�� ��Jy�3�^jY+\>��M���Ɂ�   �ً`>]���@u�M̋U�Y��
�� u�M̉�M�_3�[�k���Ë�U���|��13ŉE��E3�V3��E��EFW�E��}��M��u��M��M��M��M��M��M��M�9M$u�W����    ����3��<  �U�U��< t<	t<
t<uB��S�0�B���  �$�~Z�Hπ�wjYJ�ߋM$�	���   �	:ujY������+tHHt���|  ���jY�E� �  뤃e� jY뛍Hωu���v��M$�	���   �	:uj�<+t"<-t:�t�<C�/  <E~
,d<�!  j�Jj넍Hπ��_����M$�	���   �	:�a���:��s����U��  �u��<9�}�s
�E�*ÈG��E��B:�}�M$�	���   �	:�h���<+t�<-t��k����}� �u��u�u&��M��B:�t��<9Ճ}�s�E�*ÈG�M��B:�}��*Éu�<	�n���j�����J��M��Hπ�wj	��������+t HHt���=���j�����M��jY�Q���j�~����u���B:�t�,1<v�J�&�Hπ�v�:�뿃}  tG����+�J��M�t�HHt��у}� �E����  jX9E�v�}�|�E�O�E��E��}� ��  �Yj
YJ��
�����뾉u�3��<9 k�
���L1Ё�P  	�B:�}���Q  �M��<9�]����B:�}��Q����M��E�O�? t�E�P�u��E�P�!  �E�3҃�9U�}��E�9U�uE9U�u+E=P  �!  =�����-  �A��`�E�;���  }�عpB�E���`9Uu3�f�E�9U���  ��M�3ҋE��}���T���M�;���  k��� �  f9r��}�����M��]��U�3��E��EԉE؉E��C
��3uι�  #�#��� �  ��  ��u���f;��   f;��  ���  f;��	  ��?  f;�w3��EȉE��  3�f;�uA�E����u9u�u9u�u3�f�E���  f;�u!A�C���u9su93u�ủuȉu���  �u��}��E�   �E��U���U���~R�DĉE��C�E��E��U��� �e� �W��4;�r;�s�E�   �}� �w�tf��E��m��M��}� ����E��M��}� ����  f��~7�}܅�x+�u؋E��e����������?���  �u؉E�f���f��M����  f��yB��������E�t�E��E܋}؋U��m�������E������N�}؉E�u�9u�tf�M�� �  f9E�w�Uԁ��� �� � u4�}��u+�e� �}��u�e� ���  f9U�uf�E�A�f�E���E���Eָ�  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�M�f�EċE؉EƋE܉E�f�M��3�f�����e� H%   � ���e� �Ẽ}� �=����E��MċuƋU����/�E�   �3���  �   �3��E�   ��E�   3�3�3�3��}�E�f�f�G
�E��w�W[�M�_3�^�qd���ÍI bT�T�T0UuU�U�UVV�VwV&V��U���t��13ŉE��E�U� �  #�S�]�E��A�V#�f�}� W�]��E������E������E����?�E�   t�C-��C �u�}f��u7����   ����   3�f9M�f�����$ �Cf�C0�C 3�@�  f;���   �M3�@f��   �;�u�} t��   @uh��S3�PPPPP�g���3�f9U�t��   �u9Uu-h��;�u"9Uuh��CjP�;�������u��C�h��CjP��������u��C3��k  �ʋ�i�M  �������Ck�M��������3�f�M��عA��`�ۉE�f�U�u�}�M���  ��y�pB��`�ۉE�����  �E�T�������g  k�M����M�� �  f9r���}ĥ��Eĥ�MƉE�3ɉM��M��M�M��H
��3U��  �� �  �U��U�#�#΍4����  f;���  f;���  ���  f;���  ��?  f;�w3��u�u�u���  3�f;�uG�E����u9u�u9u�u3�f�E��  f;�uG�@���u	9pu90t�!u��u��E�   �M��U�ɉU���~U�L����M��E��E���E�� �V��ȃe� �
;�r;�s�E�   �}� �F�tf��E��m��M��}� ��E����E��M��}� ����  f��~;�E�   �u-�E�M��e��������E�E�������  �E�f���f��M����  f��yB��������E�t�E��M��u�U��m������M������H�u�M�u�9E�tf�M�� �  f9E�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�G�f�E���E���E��  f;���   3�3�f9E��E����E�I��   ��� ���M�3�;��}����M�����?  ��  f;���  �]��E�3҉U��U��U�U��U�3�#�#Ё� �  �4
�]���f;��L  f;��C  ���  f;��5  ��?  f;�wK3��E�E��9  f�E�}�f�E��E�E�E��E�f�}��Z���3�3�f9u���H%   � ���E��a���3�f;�uF�E����u9E�u9E�u	f�E���  f;�uF�E����u9E�u	9E��v����E��}��E�   �E��M���M���~K�M؉M��D��M���	�e� �ʋW��
;�r;�s�E�   �}� �_�tf��m����M��}� ����E��M��}� ����  f��~7�}���x+�E�M��e��������E����?���  �E�f���f��M����  f��yB��������E�t�E��M��}�U��m�������M������H�}�M�u�9E�tf�M�� �  f9E�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�F�f�E���E���E��  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�u�f�E��E�E�E��E�f�u��3�f�����e� H%   � ���e� �E��E�U��E��}f�t0����)3�f�� �  f9E�f�B0����$ �B�B �s�����~j_�u������?  3�f�E��E�   �E��]�M��e����؋E������M��]�E�u؅�y2�ށ��   ~(�E�]�M��m�����؋E������N�]�E���؍G�Z�]��E�����   �U��E�u��}ĥ���e��}��e���� ʋU�����֋��4	����U���ȋE���<;�r;�s�F3�;�r��s3�B����tA�Eȍ0�U�;�r;�sAM����ʍ4?�u��u��M������0������C�M��}� �u��E� �K����C���<5}�M��D�;9u	�0K;]�s�E�;]�sCf� �*؀��ˈX�D �E��M�_^3�[�[���À;0uK;�s��E�;�s�3�f�� �  f9U��@���ʀ��� �P�0�@ ����3���t@��t����t����t����t�� ��   t���˺   #�V�   t#��   t;�t;�u   �   �   �ˁ�   t��   u���^��   t   �3���t��   SVW�   ��t���t   ��t   ��t   �   ��   tǋʾ   #�t;�t;�t;�u `  � @  �    �   _#�^[��   t��   t
;�u �  Ã�@�@�  Ë�U���SVW��}�f�]�3���tjZ��t����t����t���� t����t��   �ˋ��   #ƿ   t$=   t=   t;�u����   ���   #�t��   u��   ���   �é   t��   �}�M����#�#���E;���   ���������E��m���}��]�3���tjZ��t����t����t���� t����t��   �ˋ�#�t(=   t=   t;�u��   ���   ���   ��   t��   u��   ���   ��   t��   �U��3�95tb��  ���}��]��E���yj^�   t���   t���   t���   t���   t��   �Ȼ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #ǃ�@t-�  t��@u��   ���   ���   �E��#E��#��;�u���   ����P�E������Y�]�M�3҄�yjZ��   t����   t����   t����   t���   ��t��   ��#�t$=    t= @  t;�u��   �
��   ��#σ�@t���  t��@u��   ���   ���   ��3ME�� t   �_^[������������V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� �����������U��SVWUj j h�h�u�j  ]_^[��]ËL$�A   �   t2�D$�H�3��V��U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h�hd�5    ��13�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y�hu�Q�R9Qu�   �SQ�p>�SQ�p>�L$�K�C�kUQPXY]Y[� ������������Q�L$+ȃ����Y�z  Q�L$+ȃ����Y�d  ��U��f�U��  ��f#�f;�u-�EQQ�$�����HYYtHtHt3�@]�j�jX]ø   ]��M�� �  f��u�E�� u�} t����������]��E��������D��z��������@]����%���   ]Ë�U��QQ�EV�u�E��EWV�E��Z  ���Y;�u���� 	   �ǋ��J�u�M�Q�u�P����E�;�u����t	P���Y�ϋ�����`a�����D0� ��E��U�_^��jh$�{������]܉]��E���u�I���  �.��� 	   �Ë��   ��x;Tar�!���  ���� 	   �ɦ���ы����<�`a��������L1��t�P��  Y�e� ��D0t�u�u�u�u��������E܉U���~��� 	   �~���  �]܉]��E������   �E܋U��z����u�  YË�U���  �I  ��13ŉE��EV�uW3���4�����8�����0���9}u3��  ;�u�7~���8�~���    ��������  ������S��`a������L8$�����$�����?�����t��u'�M����u��}���  �}���    聥���  �D8 tjj j V������V�>  Y����  ��D���  �k���@l3�9H�� �����P��4����3�;��`  ;�t8�?����P  ����4����� ���3���,���9E�#  ��@�����?������g  ���$���3���
��������ǃx8 t�P4�U�M��`8 j�E�P�K��P�p���Y��t:��4���+�M3�@;���  j��D���SP��  �������  C��@����jS��D���P�  ������n  3�PPj�M�Qj��D���QP�� ���C��@����t������=  j ��,���PV�E�P��$���� �4�����
  ��@�����0������8���9�,�����  ����� ��   j ��,���Pj�E�P��$���� �E��4������  ��,�����  ��0�����8����   <t<u!�33Ƀ�
������@�����D��������<t<uR��D����.  Yf;�D����I  ��8�������� t)jXP��D����  Yf;�D����  ��8�����0����E9�@���������  ����8����T4��D8��  3ɋ�D8���  ��?��� ��D�����   ��4���9M��  ��3�+�4�����H���;Ms&�CA�� �����
u��0���� @F�@F���  rՋ���H���+�j ��(���PV��H���P��$���� �4�����C  ��(����8���;��;  ��+�4���;E�l����%  ��?�����   ��4���9M�H  ��@��� ��+�4���j��H���^;MsC��Ή� �����
u�0���j[f��� �����@����@���f�Ɓ�@����  r�����H���+�j ��(���PV��H���P��$���� �4�����i  ��(����8���;��a  ��+�4���;E�G����K  ��4�����,���9M�u  ��,�����@��� +�4���j��H���^;Ms;��,�����,���΃�
uj[f���@����@���f�Ɓ�@����  r�3�VVhU  ������Q��H���+��+���P��PVh��  �t���;���   j ��(���P��+�P��5����P��$���� �4����t�(���;�������D���;�\��,���+�4�����8���;E�����?Q��(���Q�u��4����48����t��(�����D��� ��8��������D�����8��� ul��D��� t-j^9�D���u��w��� 	   ��w���0�?��D�����w��Y�1��$���� �D@t��4����8u3��$�w���    �w���  ������8���+�0���[�M�_3�^��K����jh0$�/s���]���u�kw���  �Pw��� 	   ����   ��x;Tar�Dw���  �)w��� 	   �����ҋ����<�`a�������D0��t�S��  Y�e� ��D0t�u�uS�n������E����v��� 	   ��v���  �M���E������   �E��r��Ë]S�B  YË�U���Qh   ��g��Y�M�A��t�I�A   ��I�A�A�A   �A�a �]Ë�U��E���u�Bv��� 	   3�]Å�x;Tar�'v��� 	   �����ދȃ�����`a���D��@]ø�>á@aVj^��u�   �;�}�ƣ@ajP�Wg��YY�(Q��ujV�5@a�>g��YY�(Q��ujX^�3ҹ�>��(Q��� ���� A|�j�^3ҹ�>W������`a����������t;�t��u�1�� B���>|�_3�^��
  �=�J t�p  �5(Q�?��YË�U��V�u��>;�r"���@w��+�����Q������N �  Y�
�� V���^]Ë�U��E��}��P�ʦ���E�H �  Y]ËE�� P���]Ë�U��E��>;�r=�@w�`���+�����P訥��Y]Ã� P���]Ë�U��M�E��}�`�����Q�y���Y]Ã� P���]Ë�U��E��u�8t���    ��������]Ë@]á�1��3�9Q����Ë�U���SV�u3�W�};�u;�v�E;�t�3��{�E;�t�������v��s��j^�0蒛�����V�u�M��K���E�9X��   f�E��   f;�v6;�t;�vWSV��6�����s��� *   �xs��� 8]�t�M��ap�_^[��;�t&;�w �Xs��j"^�0����8]�t��E��`p��y�����E;�t�    8]��<����E��`p��0����MQSWVj�MQS�]�p�t�;�t9]�j����M;�t�������z�P���;��s���;��k���WSV�*6�����[�����U��j �u�u�u�u������]������U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^������������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�Ë�U����ES3�VW�E�N@  ��X�X9]�E  3ɉ]���}襥��э<	���ʋU�e ��ى}����֋u����ϋ��M���U�����։0�x�H;�r;U�s�E   �} �t'�u��e �~;�r��s�E   �} �xtA�H�u�e �7;�r;�s�E   �} �XtA�HM��e� ��ɋ��������މH�M�M�M��X�1�2�u�;�r;�s�E�   �}� �t$�S3�;�r��s3�F�ډP��t
�U�B�U�P�M�U�E�} �X�P�����3�9Xu*�P��E���  ��������������P�;�t܉x�x�� �  u0�H��E���  �����������ʉ�H�x�� �  t�f�M�_^f�H
[��������������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ���U��MS3�VW;�|[;TasS��������<�`a����D0t6�<0�t0�=hDu+�tItIuSj��Sj��Sj������3���zo��� 	   �o������_^[]Ë�U��E���u�fo���  �Ko��� 	   ���]Å�x;Tar�Bo���  �'o��� 	   �����Ջ�����`a�����Dt͋]�jhP$�j���}����������4�`a�E�   3�9^u5j
辠��Y�]�9^uh�  �FP�\���u�]��F�E������0   9]�t����������`a�D8P����E��{j���3ۋ}j
耟��YË�U��E�ȃ�����`a���DP���]Ë�U��Q�=�C�u��  ��C���u���  ��j �M�Qj�MQP����t�f�E�Ë�U���SV�u3�;�t9]t8u�E;�t3�f�3�^[���u�M��E���E�9Xu�E;�t�f�8]�t�E��`p�3�@�ˍE�P�P�����YY��t}�E����   ��~%9M| 3�9]��R�uQVj	�p�ؐ���E�u�M;��   r 8^t���   8]��f����M��ap��Z����m��� *   8]�t�E��`p�����;���3�9]��P�u�E�jVj	�p�ؐ���:���뺋�U��j �u�u�u�������]�jhp$�h��3ۉ]�j覞��Y�]�j_�}�;=@a}T���(Q9�tE���@�tP��  Y���t�E��|(�(Q���� P�h��(Q�4��6��Y�(Q��G��E������	   �E��Ah���j�K���YË�U��SV�u�F�Ȁ�3ۀ�u@�  t9�FW�>+���~,WPV����YP�|�����;�u�F��y����F��N ���_�F�f �^��[]Ë�U��V�u��u	V�5   Y�/V�|���Y��t�����F @  tV�B���P�J  Y��Y��3�^]�jh�$�6g��3��}�}�j�W���Y�}�3��u�;5@a��   �(Q��98t^� �@�tVPV�G���YY3�B�U��(Q���H���t/9UuP�J���Y���t�E��9}u��tP�/���Y���u	E܉}��   F�3��u�(Q�4�V�P���YY��E������   �}�E�t�E��f���j�����Y�j����Y���������������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� 3�PPjPjh   @h������Cá�C���t���tP���Ë�U��V�uW�����u�j���    �ɑ����D�F�t8V�����V���N  V����P�~  ����y�����F��tP�4���f Y�f ��_^]�jh�$�me���M��3��u������u�i���    �O��������F@t�f �E��ye���V�<���Y�e� V�<���Y�E��E������   �ԋuV����Y�jh�$��d���]���u�"i��� 	   ����   ��x;Tar�i��� 	   �Ɛ���ڋ����<�`a�������D��t�S�����Y�e� ��Dt1S�W���YP�����u���E���e� �}� t�h���M��h��� 	   �M���E������   �E��}d��Ë]S����Y�������������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_�Ë�U��V�uWV����Y���tP�`a��u	���   u��u�@Dtj�U���j���L���YY;�tV�@���YP�����u
�����3�V����������`a����Y�D0 ��tW�g��Y����3�_^]�jh�$�c���]���u�Sg���  �8g��� 	   ����   ��x;Tar�,g���  �g��� 	   �Ԏ���ҋ����<�`a�������D0��t�S�����Y�e� ��D0tS�����Y�E���f��� 	   �M���E������   �E��b��Ë]S�:���YË�U��V�u�F��t�t�v��0���f����3�Y��F�F^]��%Đ��������h0��:��Y����̃=D uK�D��t��C�Q<P�B�Ѓ��D    �D��tV��� u��V�j������D    ^�                                                                                                                                                                                                                                                                                                                                                                                           @& P& `& v& �& �& �& �& �& �& �& �& 
' ' &' 0' H' \' l' �' �' �' �' �' �' �' ( ( 4( N( d( ~( �( �( �( �( �( �(  ) ) () D) b) v) �) �) �) �) �) �) �) �) * * &* <* N* `* p* �* �* �* �* �*          �        f����c~t        C�/u                            Gl�Q       r   � �     c:\program files\maxon\cinema 4d r12\plugins\maze trace\source\kd_tree.cpp              P�               �?c:\program files\maxon\cinema 4d r12\resource\_api\ge_dynamicarray.h    D�F p � 0� @� P�  � `� �� �� p� �� �� І �� �� �� Љ �� p� �� �� Ѝ ��   �� �� `� �� `� 0� P�     c:\program files\maxon\cinema 4d r12\plugins\maze trace\source\object\pointgenerator.cpp    Octpointgenerator   pointGenerator.tif            �?Filtering Points              @��F �3 � 0� @� P�  � `� �� �� p� �� �� І �� �� �� Љ �� p� �� �� Ѝ �� �6 �� �� `� �� `� 0� P�     c:\program files\maxon\cinema 4d r12\plugins\maze trace\source\object\tsp.cpp   Octtsp  tsp.tif error finding neighbor        �Connecting Points   Collecting Points   -DT�!��-DT�!�?-DT�!	@�������������-DT�!@�h㈵��>       @      �A      �A
ףp=
�?       �
ףp=
�?      @      @����MbP?c:\program files\maxon\cinema 4d r12\resource\_api\c4d_resource.cpp #   M_EDITOR    �Ѕ res c:\program files\maxon\cinema 4d r12\resource\_api\c4d_general.h    %s       `� � H @� c:\program files\maxon\cinema 4d r12\resource\_api\c4d_baseobject.cpp   c:\program files\maxon\cinema 4d r12\resource\_api\c4d_file.cpp c:\program files\maxon\cinema 4d r12\resource\_api\c4d_basebitmap.cpp   c:\program files\maxon\cinema 4d r12\resource\_api\c4d_libs\lib_ngon.cpp        c:\program files\maxon\cinema 4d r12\resource\_api\c4d_pmain.cpp    � 0�    c:\program files\maxon\cinema 4d r12\resource\_api\c4d_gv\ge_mtools.cpp � ��$!�p!��%��!
�          �?      �?3      3            �      0C       �       ��              e+000                  ���5�h!����?      �?            �?5�h!���>@�������             ��      �@      �        r u n t i m e   e r r o r        
     T L O S S   e r r o r  
   S I N G   e r r o r  
     D O M A I N   e r r o r  
         R 6 0 3 3  
 -   A t t e m p t   t o   u s e   M S I L   c o d e   f r o m   t h i s   a s s e m b l y   d u r i n g   n a t i v e   c o d e   i n i t i a l i z a t i o n 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .   I t   i s   m o s t   l i k e l y   t h e   r e s u l t   o f   c a l l i n g   a n   M S I L - c o m p i l e d   ( / c l r )   f u n c t i o n   f r o m   a   n a t i v e   c o n s t r u c t o r   o r   f r o m   D l l M a i n .  
     R 6 0 3 2  
 -   n o t   e n o u g h   s p a c e   f o r   l o c a l e   i n f o r m a t i o n  
     R 6 0 3 1  
 -   A t t e m p t   t o   i n i t i a l i z e   t h e   C R T   m o r e   t h a n   o n c e . 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .  
     R 6 0 3 0  
 -   C R T   n o t   i n i t i a l i z e d  
     R 6 0 2 8  
 -   u n a b l e   t o   i n i t i a l i z e   h e a p  
         R 6 0 2 7  
 -   n o t   e n o u g h   s p a c e   f o r   l o w i o   i n i t i a l i z a t i o n  
         R 6 0 2 6  
 -   n o t   e n o u g h   s p a c e   f o r   s t d i o   i n i t i a l i z a t i o n  
         R 6 0 2 5  
 -   p u r e   v i r t u a l   f u n c t i o n   c a l l  
       R 6 0 2 4  
 -   n o t   e n o u g h   s p a c e   f o r   _ o n e x i t / a t e x i t   t a b l e  
         R 6 0 1 9  
 -   u n a b l e   t o   o p e n   c o n s o l e   d e v i c e  
         R 6 0 1 8  
 -   u n e x p e c t e d   h e a p   e r r o r  
         R 6 0 1 7  
 -   u n e x p e c t e d   m u l t i t h r e a d   l o c k   e r r o r  
         R 6 0 1 6  
 -   n o t   e n o u g h   s p a c e   f o r   t h r e a d   d a t a  
   R 6 0 1 0  
 -   a b o r t ( )   h a s   b e e n   c a l l e d  
     R 6 0 0 9  
 -   n o t   e n o u g h   s p a c e   f o r   e n v i r o n m e n t  
   R 6 0 0 8  
 -   n o t   e n o u g h   s p a c e   f o r   a r g u m e n t s  
       R 6 0 0 2  
 -   f l o a t i n g   p o i n t   s u p p o r t   n o t   l o a d e d  
            ��   P�	   ��
   ��   X�   ��   ��   X�   �   ��   (�   ��   h�   (�   `�    ��!   �x   �y   Șz   ���   ���   ��M i c r o s o f t   V i s u a l   C + +   R u n t i m e   L i b r a r y     
 
     . . .   < p r o g r a m   n a m e   u n k n o w n >     R u n t i m e   E r r o r ! 
 
 P r o g r a m :     K E R N E L 3 2 . D L L     FlsFree FlsSetValue FlsGetValue FlsAlloc    CorExitProcess  m s c o r e e . d l l     �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       � �       � �          	   �                    8C      8CX������< 1�
�"�?'���;�< ï&�b�?�,kg��< !J���?ĂeT1��< �1y"�?�z���< �F#�?V���a�< $�
lc�?���x��< �nu���?c�v5��< ����?0��N�< �ߢ�#�?	��"$�< b�md�?�g�Q��< |a7��?�麏��< a��c�?0H_��< �А$�?]U ?�< 8�U�d�?|}}�?�< 5�盧?~+����<  �?)0>�B��< �'HR%�?���I&�< ^:ȅe�?>!ʎ��< sl����?e�cb~q�< �ۧ��?r���ʀ�< F�(&�?Z��n��< '��`f�?4�7j��< ��㚦�?+i��	U�< �oX��?F��.K;�< ��.'�?Yh�ŉ�< 4lkQg�?�;+�U��< 3���?�М	m8�< ��&��?����< �S�(�?Y�=�t< :@�Xh�?,�n@4`�< ��$���?�����< �n��?��9�ܮ�< � �-)�?\�����< �Řwi�?���=�< R�%é�?�f�@��< *�B�?a���w��< G��^*�?�m(�<��< �2;�j�?��P�E�< ����?<�/����< :�T�?Ft����< ͩ+�?N�ibzP�< ��� l�?��  %X�< aY��?]@�_}�< �nL��?����G	�< �1-�?a���(�< U�lm�?iT	�?��< �*̭�?V��*���< w7H-�?��X[F�< �+�.�?X� kn�< E���n�?�T�(�+�< ��U[��?։���< '���?ju!4���< ��-0�?������< Q̙p�?�冿��< �����?���{��< qw�?_W����< �C�1�?'����< I��\r�?��D�c< s�>Ҳ�?������< w*�I�?���n'$�< �2�3�?z���7�< [��>t�?V-Ai��< �����?`�DTb�< �;��?S��.��< TR�*�?)�R���< 2���k�?,�%�ً�< r����?SC?
�< H����?Zxg�f��< �`/-�?����#�< މ7�m�?�w���< 悆a��?_"�C���< lX^��?���@��< �{Х/�?$�8�^�< ]h�Np�?b�X*��< �����?�}�_Ͼ< ��s���?��p�t�< �h�f2�?��$�V�< �4{#s�?U���g
�< ����?��w���< J.����?I�Z��< *�Ow5�?��.@��< ��FHv�?N	����< �!���?�j����< �v(���?��z�"�< i�6�8�? �?!���< <���y�?G��o��< �魺�?�xeF���< �豟��?�G��T��< ��1�<�?V�	ڀ�< ��{�}�?���0���< �����?���a@��< ﶠ��?�0����< ��̯@�?��1�< �3�ā�?��.aU�< !�E���?�I�����< ����?���	���< �j�)E�?O�����< I�W��?W�0�e)�< ��u���?����
T�< �˛��?����?��< �X	J�?!PO79�< �/�Q��?�;�X��< J]���?V:e:���< �Q���?�Wm��`�< b;�SO�?4Td'��< 
Xw���?ЀY��< �L"��?d��ݩS�< _}?��?�T�x�< �[bU�?�\�z#��< ^ɍ��?1����< �N���?�wa���< �����?���N9�< a�X;[�?���Y']�< @ٜ̓�?���E�< VOu��?!S�ÀX�< b- �?C�:���< �|�a�?B�<��$�< �{ɟ��?+X�UG�< m�e��?>Uۊ�< �o]2'�?�� I��< Р�i�?G�����< ��o��? ��Ιn�< 9�[���?�	�|�^�< ����.�?�>oj��< .�_�p�?1S���< �X����?����l�< �~���?o.x���< %3d�?����{ = 4 ��L�?�V!�= b�#��?��@g	= a��?G��z	= �]ư�?���6�= o�JV�?J�� �b= '4��?/��t�>�< w���?a�`����< �_��?a�	�e= ��F``�?/�f	= #&��?�5SmT4�< W�� ��?R�z��<  ъ�(�?���vY�< ���k�?p�Y�.= �y���?�8�'���< Ku�C��?j��<{= 2�<�5�?��ýd	= ��x�?�"a��= @�ic��?�%�[�9= �����?kR�F��< �6D�C�?ş
ܬ_�< 5��Z��?ȡ�k*= ���3��?�*+xi(�< �G�&�?��r
ly= :��3S�?z
�j�< �[��?��'����< ;!���?h����= �<��?���:��< ��sd�?��3�= �?	��?{�!m�B�< <>����?�*�2 = ����2�?cM�yoG= V��sw�?8K��$�< ��}��?C�l���< Ϲ���?�-��< '���F�?ɕ���{�< �$�R��?܊�)B��< �#���?������< ��c�?? ��~��< ���F]�?���&��= �		/��?94��E�< ?T9��?9*��)�< l?�e/�?�B6�!F= u0w�u�?�M�떐= �k`(��?������< 4�=��?Kp��= G"�zI�?$�}Tw5�< �[��?ߪ��b�< �Ka��?aF7�= Vj��?�T��y�< R߂�e�?M]-��e�< $�[��?3����< Ễ���?��QZo�= n��<�?1-
I�x�< f�	���?I��]�= ��O���?���x�= �#$�?�nz��= �) �]�?����h��< �'�7��?y]h�= �Yg��?�S�c�< b}��?��$ګ= ;�ђ@�?OD���)= ���=e�?:Q�]D\�< ��� ��?FnH�AY�< "�ۮ�?�)Bp�= )R�Q��?��{���< �L��0�?�U��< d�N{�?���c�1= f��k��?iO��)= ��m��?�
��R = l[��]�?�$Ŝi= w/�d��?���C�= �(�O��?u��1��= ��/�D�? �&= �� ���?i�C1]�< Ei��?X�=g��< P�~0�?Y;���=  ]��?���m��< �����?�A�8�y�< �7�l �?S6���= =.�q�?+`���= �����?���%!5= �o�h�?�y���= i�Q�i�?v�7���= �Խ�?dDR޸;= nl���?b*t#�= x�A@h�?�����= ZmI���?�oP�@= ��Y��?��Ͽ	= �n�?u�И?�= %�k��?ZEM-'^= DT!�?:Z��n== ��0|�?�O���= ���*��?m}I�{= �eP5�?+�}ZI= �Q����?�^oc;�< '��?
u�/r��< ���S�?�i���1= �q���?/����= {�ss�?VV&�= �#�k~�?[��	�< �����?vB���< 6��#M�?��!��< 
��?q_�w#�< ����"�?ұ��R��< �����?k=�C= �B� �?��_���< u���r�?�y���= Dw�b��?�(,xn�< <"Q/�?���q�q)= �o\l�?�)���T&=  7a��?��L�< �?|6��?�������?#�DZ9��?������?��/�.��?>6)}���?, �,��?��؏��?M�����?��x%q��?�� ����?/x�bJ��?Ȉb����?�uÏ��?(Z����?��t����?{}�2F��?�������?_�2��?>�T�^��?�u	���?�����?4t��d��?��Z���?(�	��?WI�Y��?�d���?�{�����?|��:��?�S9���?���s���?���
��?����K��??�����?l�.���?�Z�3��?��;E<��?�fSOs��?�J�Q���?�z�L���?�@��?{yK+;��?ãjh��?��F���?-(�����?�n�����?@��F��?����)��?�P�J��?C��Si��?�^����?�B����?i|e���?�������?�� ���?�a�k���?c����?X�!��?89�l!��?fh�+��?��3��?)Ao
:��?�1(>��?2:@��?>�?@@��?"I�r���?6��4���?�@Û��?����?765@Z��?�&+-��?w�'����?��Q���?�Gp�t��?�2�&��?X��9Ш�?B�q��?/�?�
��?v�ɛ��?��Mj$��?�3����?�s����?b里��?V�����?%S��?V��ѩ��?ߖ%@���?�U>��?2�,|��?�ܜm���?V��kށ�?9�?�I�@|�?��P3y�?�?}>v�?��H|As�?#�<p�?_0.m�?t���j�?���f�?�����c�?�3)�`�?��i]�?�� F)Z�?�2V�V�?��f\�S�?B?}4P�?���V�L�?{�fI�?uS�E�?|�ǩuB�?1�<��>�?�(��b;�?�탿�7�?�]o�-4�?P�h�0�?�H�,�?�:5�)�?Iٓ\%�?f,��!�?갸%��?N���?$�k��?�oay�?*���?��?Y
�?���$�?�?�(�?���a���?�9y����?99R��?%��R���?F�����?��@�I��?j �T��?�0<��?2j���?�p�~���?,�L��?@�_�o��?7�����?�'�����?�VG��?�D<xZu�?`\@��j�?)]G�q`�?L�c�U�?�Jup�J�?CY���?�?� X7�4�?�T��)�?KB	�0�?&D��?lU����?�E0d��?KYC ��?�:����?@М����?��L���?#�e�m��?-Fգ��?�DT����?�W�㗖�?*�MU��?�z��{�?�l�Un�?
Q-��`�?>�ұR�?V�D��D�?oW�sg6�?U��J(�?>��t�?2̄λ
�?�1_����?$*2���?[��ێ��?N��)��?���V���?l$G~ٮ�?��+6��?�tF4؎�?��,�~�?����"n�?<�փ]�?|ߠ�L�?l6���;�?6*��*�?�|�59�?��:��?H�K����?s7��?��I-���?�$z����?�9\���?��>|.~�?�-��W�?�^\sY0�?:Rp�7�?m�bzA��?G�4's��?I�y�Ȋ�?%��=_�?�C\�2�?�O��u�?�m��.��?�M����?���n�w�?KK�'�F�?��l^�?:��" ��?��Ѭ�?��}6lw�?�:�@�? 7Z8>	�?$�� f��?e')lW��?zD@	[�?���jq�?�P J���?F���<��?�Q'J�`�?x��e_�?* Aӱ��?�"�Sr��?xw��N�?k��$��?
�S/���?��yx|o�?P�6 d!�?ZyrI��?�����?��Ӳ�*�?
T�����?���!�z�?��{��?��0�V��?�8I�^�?��A;��?���wC��?�JG7�&�?�'un�?���)��?m���y��?������?��|�ȕ�?,"��Q��?�/��b�?PV3� 2�?�S����?p����?V�a��"�?�Tl��?Pq�j��?��Y��?p�,�?�l"։�?cY�����?\3&��<-DT�!�?       �           �����   �����    ���UUUUUU�?333333�?�m۶mۦ?颋.��?333333�?�q�q�?UUUUUU�?O��N�đ?�m۶mۦ?$rxxx��?�������?�������     ���      �?       �9��B.�@  ׽2b      �              8C      8CX������< 1�
�"�?'���;�< ï&�b�?�,kg��< !J���?ĂeT1��< �1y"�?�z���< �F#�?V���a�< $�
lc�?���x��< �nu���?c�v5��< ����?0��N�< �ߢ�#�?	��"$�< b�md�?�g�Q��< |a7��?�麏��< a��c�?0H_��< �А$�?]U ?�< 8�U�d�?|}}�?�< 5�盧?~+����<  �?)0>�B��< �'HR%�?���I&�< ^:ȅe�?>!ʎ��< sl����?e�cb~q�< �ۧ��?r���ʀ�< F�(&�?Z��n��< '��`f�?4�7j��< ��㚦�?+i��	U�< �oX��?F��.K;�< ��.'�?Yh�ŉ�< 4lkQg�?�;+�U��< 3���?�М	m8�< ��&��?����< �S�(�?Y�=�t< :@�Xh�?,�n@4`�< ��$���?�����< �n��?��9�ܮ�< � �-)�?\�����< �Řwi�?���=�< R�%é�?�f�@��< *�B�?a���w��< G��^*�?�m(�<��< �2;�j�?��P�E�< ����?<�/����< :�T�?Ft����< ͩ+�?N�ibzP�< ��� l�?��  %X�< aY��?]@�_}�< �nL��?����G	�< �1-�?a���(�< U�lm�?iT	�?��< �*̭�?V��*���< w7H-�?��X[F�< �+�.�?X� kn�< E���n�?�T�(�+�< ��U[��?։���< '���?ju!4���< ��-0�?������< Q̙p�?�冿��< �����?���{��< qw�?_W����< �C�1�?'����< I��\r�?��D�c< s�>Ҳ�?������< w*�I�?���n'$�< �2�3�?z���7�< [��>t�?V-Ai��< �����?`�DTb�< �;��?S��.��< TR�*�?)�R���< 2���k�?,�%�ً�< r����?SC?
�< H����?Zxg�f��< �`/-�?����#�< މ7�m�?�w���< 悆a��?_"�C���< lX^��?���@��< �{Х/�?$�8�^�< ]h�Np�?b�X*��< �����?�}�_Ͼ< ��s���?��p�t�< �h�f2�?��$�V�< �4{#s�?U���g
�< ����?��w���< J.����?I�Z��< *�Ow5�?��.@��< ��FHv�?N	����< �!���?�j����< �v(���?��z�"�< i�6�8�? �?!���< <���y�?G��o��< �魺�?�xeF���< �豟��?�G��T��< ��1�<�?V�	ڀ�< ��{�}�?���0���< �����?���a@��< ﶠ��?�0����< ��̯@�?��1�< �3�ā�?��.aU�< !�E���?�I�����< ����?���	���< �j�)E�?O�����< I�W��?W�0�e)�< ��u���?����
T�< �˛��?����?��< �X	J�?!PO79�< �/�Q��?�;�X��< J]���?V:e:���< �Q���?�Wm��`�< b;�SO�?4Td'��< 
Xw���?ЀY��< �L"��?d��ݩS�< _}?��?�T�x�< �[bU�?�\�z#��< ^ɍ��?1����< �N���?�wa���< �����?���N9�< a�X;[�?���Y']�< @ٜ̓�?���E�< VOu��?!S�ÀX�< b- �?C�:���< �|�a�?B�<��$�< �{ɟ��?+X�UG�< m�e��?>Uۊ�< �o]2'�?�� I��< Р�i�?G�����< ��o��? ��Ιn�< 9�[���?�	�|�^�< ����.�?�>oj��< .�_�p�?1S���< �X����?����l�< �~���?o.x���< %3d�?����{ = 4 ��L�?�V!�= b�#��?��@g	= a��?G��z	= �]ư�?���6�= o�JV�?J�� �b= '4��?/��t�>�< w���?a�`����< �_��?a�	�e= ��F``�?/�f	= #&��?�5SmT4�< W�� ��?R�z��<  ъ�(�?���vY�< ���k�?p�Y�.= �y���?�8�'���< Ku�C��?j��<{= 2�<�5�?��ýd	= ��x�?�"a��= @�ic��?�%�[�9= �����?kR�F��< �6D�C�?ş
ܬ_�< 5��Z��?ȡ�k*= ���3��?�*+xi(�< �G�&�?��r
ly= :��3S�?z
�j�< �[��?��'����< ;!���?h����= �<��?���:��< ��sd�?��3�= �?	��?{�!m�B�< <>����?�*�2 = ����2�?cM�yoG= V��sw�?8K��$�< ��}��?C�l���< Ϲ���?�-��< '���F�?ɕ���{�< �$�R��?܊�)B��< �#���?������< ��c�?? ��~��< ���F]�?���&��= �		/��?94��E�< ?T9��?9*��)�< l?�e/�?�B6�!F= u0w�u�?�M�떐= �k`(��?������< 4�=��?Kp��= G"�zI�?$�}Tw5�< �[��?ߪ��b�< �Ka��?aF7�= Vj��?�T��y�< R߂�e�?M]-��e�< $�[��?3����< Ễ���?��QZo�= n��<�?1-
I�x�< f�	���?I��]�= ��O���?���x�= �#$�?�nz��= �) �]�?����h��< �'�7��?y]h�= �Yg��?�S�c�< b}��?��$ګ= ;�ђ@�?OD���)= ���=e�?:Q�]D\�< ��� ��?FnH�AY�< "�ۮ�?�)Bp�= )R�Q��?��{���< �L��0�?�U��< d�N{�?���c�1= f��k��?iO��)= ��m��?�
��R = l[��]�?�$Ŝi= w/�d��?���C�= �(�O��?u��1��= ��/�D�? �&= �� ���?i�C1]�< Ei��?X�=g��< P�~0�?Y;���=  ]��?���m��< �����?�A�8�y�< �7�l �?S6���= =.�q�?+`���= �����?���%!5= �o�h�?�y���= i�Q�i�?v�7���= �Խ�?dDR޸;= nl���?b*t#�= x�A@h�?�����= ZmI���?�oP�@= ��Y��?��Ͽ	= �n�?u�И?�= %�k��?ZEM-'^= DT!�?:Z��n== ��0|�?�O���= ���*��?m}I�{= �eP5�?+�}ZI= �Q����?�^oc;�< '��?
u�/r��< ���S�?�i���1= �q���?/����= {�ss�?VV&�= �#�k~�?[��	�< �����?vB���< 6��#M�?��!��< 
��?q_�w#�< ����"�?ұ��R��< �����?k=�C= �B� �?��_���< u���r�?�y���= Dw�b��?�(,xn�< <"Q/�?���q�q)= �o\l�?�)���T&=  7a��?��L�< �?|6��?�������?#�DZ9��?������?��/�.��?>6)}���?, �,��?��؏��?M�����?��x%q��?�� ����?/x�bJ��?Ȉb����?�uÏ��?(Z����?��t����?{}�2F��?�������?_�2��?>�T�^��?�u	���?�����?4t��d��?��Z���?(�	��?WI�Y��?�d���?�{�����?|��:��?�S9���?���s���?���
��?����K��??�����?l�.���?�Z�3��?��;E<��?�fSOs��?�J�Q���?�z�L���?�@��?{yK+;��?ãjh��?��F���?-(�����?�n�����?@��F��?����)��?�P�J��?C��Si��?�^����?�B����?i|e���?�������?�� ���?�a�k���?c����?X�!��?89�l!��?fh�+��?��3��?)Ao
:��?�1(>��?2:@��?>�?@@��?"I�r���?6��4���?�@Û��?����?765@Z��?�&+-��?w�'����?��Q���?�Gp�t��?�2�&��?X��9Ш�?B�q��?/�?�
��?v�ɛ��?��Mj$��?�3����?�s����?b里��?V�����?%S��?V��ѩ��?ߖ%@���?�U>��?2�,|��?�ܜm���?V��kށ�?9�?�I�@|�?��P3y�?�?}>v�?��H|As�?#�<p�?_0.m�?t���j�?���f�?�����c�?�3)�`�?��i]�?�� F)Z�?�2V�V�?��f\�S�?B?}4P�?���V�L�?{�fI�?uS�E�?|�ǩuB�?1�<��>�?�(��b;�?�탿�7�?�]o�-4�?P�h�0�?�H�,�?�:5�)�?Iٓ\%�?f,��!�?갸%��?N���?$�k��?�oay�?*���?��?Y
�?���$�?�?�(�?���a���?�9y����?99R��?%��R���?F�����?��@�I��?j �T��?�0<��?2j���?�p�~���?,�L��?@�_�o��?7�����?�'�����?�VG��?�D<xZu�?`\@��j�?)]G�q`�?L�c�U�?�Jup�J�?CY���?�?� X7�4�?�T��)�?KB	�0�?&D��?lU����?�E0d��?KYC ��?�:����?@М����?��L���?#�e�m��?-Fգ��?�DT����?�W�㗖�?*�MU��?�z��{�?�l�Un�?
Q-��`�?>�ұR�?V�D��D�?oW�sg6�?U��J(�?>��t�?2̄λ
�?�1_����?$*2���?[��ێ��?N��)��?���V���?l$G~ٮ�?��+6��?�tF4؎�?��,�~�?����"n�?<�փ]�?|ߠ�L�?l6���;�?6*��*�?�|�59�?��:��?H�K����?s7��?��I-���?�$z����?�9\���?��>|.~�?�-��W�?�^\sY0�?:Rp�7�?m�bzA��?G�4's��?I�y�Ȋ�?%��=_�?�C\�2�?�O��u�?�m��.��?�M����?���n�w�?KK�'�F�?��l^�?:��" ��?��Ѭ�?��}6lw�?�:�@�? 7Z8>	�?$�� f��?e')lW��?zD@	[�?���jq�?�P J���?F���<��?�Q'J�`�?x��e_�?* Aӱ��?�"�Sr��?xw��N�?k��$��?
�S/���?��yx|o�?P�6 d!�?ZyrI��?�����?��Ӳ�*�?
T�����?���!�z�?��{��?��0�V��?�8I�^�?��A;��?���wC��?�JG7�&�?�'un�?���)��?m���y��?������?��|�ȕ�?,"��Q��?�/��b�?PV3� 2�?�S����?p����?V�a��"�?�Tl��?Pq�j��?��Y��?p�,�?�l"։�?cY�����?\3&��<-DT�!�?\3&���-DT�!	�\3&��<-DT�!	@       �           �����   �����    ���                UUUUUUſ333333���m۶mۦ�颋.��?333333�?�q�q�?UUUUUU�?O��N�đ?�m۶mۦ?$rxxx��?�������?�������     ���      �?      �?       �9��B.�@  ׽2b      �              �7                              �?1mm.�s�,�)���?   �'>�      �?�i����i<���?   �mb�      �?Z"�������.��?   ���u�      �?ϕk��|��c����}�?   ��,g�      �?y�sh:��;�8]+�?    �^<      �?ty�[g�ſ�h�9;��?    �%�<      �?���S�Ϳ�	%�L�?    jh<      �?2���y��?�;f���?    4݋�      �?Xw$��3�?Ak���?    �ł�      �?��暳s�?��)f��?   �0�9<      �?N��,J������8�?   ���v�      �?uZEeu��F�2�k��?    �Wt<      �?-��v1��?�-�VA��?   �`�<      �?�gY���\�ϗb�?    bu<      �?P/Ye���&%ѣ���?   @�}��      �?              �?                P/Ye��?&%ѣ���?   @�}��      ���gY�?�\�ϗb�?    bu<      п-��v1����-�VA��?   �`�<      пuZEeu�?F�2�k��?    �Wt<      �N��,J�?����8�?   ���v�      ࿇�暳s����)f��?   �0�9<      �Xw$��3��Ak���?    �ł�      �2���y�ʿ�;f���?    4݋�      ����S��?�	%�L�?    jh<      �ty�[g��?�h�9;��?    �%�<      �y�sh:�?;�8]+�?    �^<      �ϕk��|�?c����}�?   ��,g�      �Z"����?��.��?   ���u�      ��i��?�i<���?   �mb�      �1mm.�s?,�)���?   �'>�      �                              �1mm.�s?,�)����   �'><      ��i��?�i<��ȿ   �mb<      �Z"����?��.�ҿ   ���u<      �ϕk��|�?c����}ؿ   ��,g<      �y�sh:�?;�8]+޿    �^�      �ty�[g��?�h�9;��    �%��      ����S��?�	%�L�    jh�      �2���y�ʿ�;f���    4݋<      �Xw$��3��Ak���    �ł<      ࿇�暳s����)f��   �0�9�      �N��,J�?����8�   ���v<      �uZEeu�?F�2�k��    �Wt�      �-��v1����-�VA��   �`��      п�gY�?�\�ϗb�    bu�      пP/Ye��?&%ѣ���   @�}�<      ��              �                P/Ye���&%ѣ���   @�}�<      �?�gY���\�ϗb�    bu�      �?-��v1��?�-�VA��   �`��      �?uZEeu��F�2�k��    �Wt�      �?N��,J������8�   ���v<      �?��暳s�?��)f��   �0�9�      �?Xw$��3�?Ak���    �ł<      �?2���y��?�;f���    4݋<      �?���S�Ϳ�	%�L�    jh�      �?ty�[g�ſ�h�9;��    �%��      �?y�sh:��;�8]+޿    �^�      �?ϕk��|��c����}ؿ   ��,g<      �?Z"�������.�ҿ   ���u<      �?�i����i<��ȿ   �mb<      �?1mm.�s�,�)����   �'><      �?UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      ��������                                      �?1mm.�s�,�)���?   �'>�      �?�i����i<���?   �mb�      �?Z"�������.��?   ���u�      �?ϕk��|��c����}�?   ��,g�      �?y�sh:��;�8]+�?    �^<      �?ty�[g�ſ�h�9;��?    �%�<      �?���S�Ϳ�	%�L�?    jh<      �?2���y��?�;f���?    4݋�      �?Xw$��3�?Ak���?    �ł�      �?��暳s�?��)f��?   �0�9<      �?N��,J������8�?   ���v�      �?uZEeu��F�2�k��?    �Wt<      �?-��v1��?�-�VA��?   �`�<      �?�gY���\�ϗb�?    bu<      �?P/Ye���&%ѣ���?   @�}��      �?              �?                P/Ye��?&%ѣ���?   @�}��      ���gY�?�\�ϗb�?    bu<      п-��v1����-�VA��?   �`�<      пuZEeu�?F�2�k��?    �Wt<      �N��,J�?����8�?   ���v�      ࿇�暳s����)f��?   �0�9<      �Xw$��3��Ak���?    �ł�      �2���y�ʿ�;f���?    4݋�      ����S��?�	%�L�?    jh<      �ty�[g��?�h�9;��?    �%�<      �y�sh:�?;�8]+�?    �^<      �ϕk��|�?c����}�?   ��,g�      �Z"����?��.��?   ���u�      ��i��?�i<���?   �mb�      �1mm.�s?,�)���?   �'>�      �                              �1mm.�s?,�)����   �'><      ��i��?�i<��ȿ   �mb<      �Z"����?��.�ҿ   ���u<      �ϕk��|�?c����}ؿ   ��,g<      �y�sh:�?;�8]+޿    �^�      �ty�[g��?�h�9;��    �%��      ����S��?�	%�L�    jh�      �2���y�ʿ�;f���    4݋<      �Xw$��3��Ak���    �ł<      ࿇�暳s����)f��   �0�9�      �N��,J�?����8�   ���v<      �uZEeu�?F�2�k��    �Wt�      �-��v1����-�VA��   �`��      п�gY�?�\�ϗb�    bu�      пP/Ye��?&%ѣ���   @�}�<      ��              �                P/Ye���&%ѣ���   @�}�<      �?�gY���\�ϗb�    bu�      �?-��v1��?�-�VA��   �`��      �?uZEeu��F�2�k��    �Wt�      �?N��,J������8�   ���v<      �?��暳s�?��)f��   �0�9�      �?Xw$��3�?Ak���    �ł<      �?2���y��?�;f���    4݋<      �?���S�Ϳ�	%�L�    jh�      �?ty�[g�ſ�h�9;��    �%��      �?y�sh:��;�8]+޿    �^�      �?ϕk��|��c����}ؿ   ��,g<      �?Z"�������.�ҿ   ���u<      �?�i����i<��ȿ   �mb<      �?1mm.�s�,�)����   �'><      �?UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      �      �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��tan cos sin modf    floor   ceil    atan    exp10   acos    asin    log log10   exp pow       �      ���������������-DT�!�?-DT�!��RUUUUU�?        v�F�$I�?������ɿ��3Y�E�?#Y��q���n����?��;
9��� ��/I�?hK����d��?81�U����H!G�?��#�$�����0|f?�K�RVn���TUUUU�?        ~I�$I�?g����ɿHB�;E�?����q���{雮?�x��֚��                   �      �?       @       @      �?      �?      @>��1|�MC              ������ ������ ������B������B  �����  ����� 8��B.�?0gǓW�.=        ����������������              �?      �?                      0C      0C      ��      �     �     �U�	�I�? ���Ͽu}�M�Uſ�UUUUU�?Sz�����?     �      �?      �?     ��?     ��?     �?     �?     ��?     ��?     �?     �?     ��?     ��?     B�?     B�?     ��?     ��?     r�?     r�?     �?     �?     ��?     ��?     N�?     N�?     ��?     ��?     ��?     ��?     B�?     B�?     ��?     ��?     ��?     ��?     H�?     H�?     ��?     ��?     ��?     ��?     b�?     b�?     �?     �?     ��?     ��?     ��?     ��?     F�?     F�?     �?     �?     ��?     ��?     ��?     ��?     B�?     B�?     �?     �?     ��?     ��?     ��?     ��?     V�?     V�?     �?     �?     ��?     ��?     ��?     ��?     z�?     z�?     F�?     F�?     �?     �?     ��?     ��?     ��?     ��?     ��?     ��?     R�?     R�?     $�?     $�?     ��?     ��?     ��?     ��?     ��?     ��?     t�?     t�?     J�?     J�?      �?      �?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     \�?     \�?     6�?     6�?     �?     �?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     b�?     b�?     B�?     B�?      �?      �?      �?      �?                  <����?N~�'��<  x�z�?��'�*$=  �#�f�?�$/��= @�0�?@A�S��1= �c�E�?�Pa�B== `�R�?Dj0Q:W$= ��>m��?��Lyc>= �*p%�?���?C;0= ��|���?�Ix�"�<= ``ә�?��y M== �or�O�?��+C��== ��v��?�����R1= PQ	��?��Ӏb= @��P�?�5M[g?= �V���?d+��[7= ������?n��B�>=  kz�*�?�w�#8= 0�nط�?C�#�7= �{���?Di�00= �ˮf�?�j -= x���)�?���}z�=  ����?��0$= H�V��?����o�= X��a�?��;�M_8= @��?�����5= ����?�^���@'= �L$��?��/r(= � <�?�vT�� 3= ��?���?��Cg��?= 0��Ә�?W/f�1= `(J�?Dk����0= h��#��?@� �6= �۫���?��_��= �|�D�?�&�?4j<= '����?Q���n�&= �ַ��?�l����= �Ð6�?�DX�,4= �����?��-Q�2= �xb�t�?�W��E��< �.l�?��7�w�,= ���Ȭ�?l�>= �ɥ�%�?��Nl,"= �@\r�?�?� t�8= 85�R��?ӇӜ��= L.��	�?�>)g�= Ը�3U�?�Ӱ��== �����?h���Xg+= �og���?�����X= ��ذ0�?{fHn�= <��w�?y�5s3R6= ��)��?��a8��< O4W�?4�bV�0= ����L�?�4���@= ���@��?�X��ۓ4= Tk���?>�_��(=  ����?�*��o= �@�[c�?�����,= $4b��?d����O"= lx���?#60���8= ě&m*�?ɉ�h"0= �בl�?�n6ѯ{�< 9[P��?�ce�zb�< $����?�F�8"= 8��B.�?0gǓW�.=       ��       ���ܧ׹�fq�@      ��@�6C����?      �?exp          ����  L`LH H : m m : s s     d d d d ,   M M M M   d d ,   y y y y   M M / d d / y y     P M     A M     D e c e m b e r     N o v e m b e r     O c t o b e r   S e p t e m b e r   A u g u s t     J u l y     J u n e     A p r i l   M a r c h   F e b r u a r y     J a n u a r y   D e c   N o v   O c t   S e p   A u g   J u l   J u n   M a y   A p r   M a r   F e b   J a n   S a t u r d a y     F r i d a y     T h u r s d a y     W e d n e s d a y   T u e s d a y   M o n d a y     S u n d a y     S a t   F r i   T h u   W e d   T u e   M o n   S u n   HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun  Complete Object Locator'    Class Hierarchy Descriptor'     Base Class Array'   Base Class Descriptor at (  Type Descriptor'   `local static thread guard' `managed vector copy constructor iterator'  `vector vbase copy constructor iterator'    `vector copy constructor iterator'  `dynamic atexit destructor for '    `dynamic initializer for '  `eh vector vbase copy constructor iterator' `eh vector copy constructor iterator'   `managed vector destructor iterator'    `managed vector constructor iterator'   `placement delete[] closure'    `placement delete closure'  `omni callsig'   delete[]    new[]  `local vftable constructor closure' `local vftable' `RTTI   `EH `udt returning' `copy constructor closure'  `eh vector vbase constructor iterator'  `eh vector destructor iterator' `eh vector constructor iterator'    `virtual displacement map'  `vector vbase constructor iterator' `vector destructor iterator'    `vector constructor iterator'   `scalar deleting destructor'    `default constructor closure'   `vector deleting destructor'    `vbase destructor'  `string'    `local static guard'    `typeof'    `vcall' `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ~   ()  ,   >=  >   <=  <   %   /   ->* &   +   -   --  ++  *   ->  operator    []  !=  ==  !   <<  >>  =    delete  new    __unaligned __restrict  __ptr64 __eabi  __clrcall   __fastcall  __thiscall  __stdcall   __pascal    __cdecl __based(    <�4�(��������������ӑ��������������������������������|�x�t�p�l�h�d�`�\�X�T�P�L�H�D�@�<�8�4�0�,�(�$� ����������������x�X�8����������l�P�@�<�4�$� �����������x�P�(���������l�@�$�ӑ���������GetProcessWindowStation GetUserObjectInformationW   GetLastActivePopup  GetActiveWindow MessageBoxW U S E R 3 2 . D L L     _nextafter  _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   fabs    sqrt    atan2   tanh    cosh    sinh       �U��?�wB%�K�=      �?   �[��?(�6N�g�=      �?   $�?V�`t� >      �?   ��տ?��2n{a>      �?   ����?��M��=      �?   H{��?{4�r>      �?   Pא�?"�"�>      �?   �u[�?��*��>      �?   ����?G�0��_(>      �?   4wb�?��i^^?(>      �?   ��0�?p3���>      �?   @��?F��M>      �?   8M��?�B�V��>      �?   ��d�?}B��a.>      �?   ȴ�?d�����>      �?   g��?�ߊ��>      �?   �@�?�f\���*>      �?   �~e�?�-��f>      �?   �]%�?D	�G��?>      �?   ���?�\����>>      �?   X���?�1��#>      �?   �E�?��h��>      �?   �?��?�ⳇ��>      �?   ����?�$	�49>      �?   x�8�?k���0H<>      �?   ����?r��ش8>      �?   8fm�?�"m>">      �?   ħ �?[��<c�'>      �?   �k��?"���%>      �?   ���?݉@fR�8>      �?   ����?��T���:>      �?   T�!�?3&�F>      �?   � ��?<����[#>     ��?   �%�?�Y:/(A6>      �?   ����?��N��2>     ��?   8O�?�r�!'	>      �?   ��r�?���8{K>     ��?   �p��?9��l�9$>      �?   �
G�?�aj	�i9>     ��?   T|��?'\�|#<>      �?   $��?�}�dj�#>     ��?   �Wn�?׈MVx:>      �?   ,���?1�8o,>     ��?   D�$�?	c�/�
>      �?   @ |�?��x7|�1>     ��?   |���?��9>      �?   p #�?�IA��u=>     ��?   �s�?�x ٴ4>      �?   p���?edf�&�.>     ��?   ,�?��f���A>      �?   h�*�?v����2>     ��?   $gN�?RE\��K>      �?   �q�?'^��IE>     ��?   DΒ�?��&a��H>      �?   L���?�&KrQF>     ��?   ,���?�#/�'�>      �?   إ��?]X�c�?>     ��?    ��?�Ԯ}�>      �?   �e.�?�IdW�A>     ��?   �K�?���ΐ?>      �?   Xg�?��4*�A>     ��?   _��?�[�ǆJ>      �?   ���?1���0H>     ��?   ���?�hc#�]G>       @   ,*��?�Q�x
�F>     @ @   p���?ek�R�.N>     � @   �� �?�Ӿ�n@>     � @   �b�?�����O>      @   $Q/�?CJ���O>     @@   ��E�?������G>     �@   �[�?�3E�{A>     �@   T�p�?�SfI�S:>      @   X΅�?B6)�1�<>     @@   �3��?>ځ���7>     �@   $��?s(��N>     �@   @���?V�
6�f=>      @   (���?��{��>     @@   (W��?��-�Jg >     �@   ����?��"a�PK>     �@   xm�?,S��ڤ6>      @   ���?�6��hb">     @@    �-�?�k,�<>     �@   X�>�?�0����=>     �@   �O�?�׀IX�H>      @   �-_�?���
@>     @@   ��n�?���2E>     �@   �P~�?�=�ő�8>     �@   lj��?�[j&,>      @   L7��?��x��82>     @@   ����?c�#V�B>     �@   0��?7ڨ.�Y>     �@   P���?�[�p&>      @   ؔ��?h4�M��A>     @@   � ��?E�p�l E>     �@   �+��?�o�$�E>     �@   h��?\���*�K>      @   ���?-�?��B>     @@   P8�?�(l�|�@>     �@   �p!�?u���@�J>     �@   @p-�?�V��1>      	@   �89�?����5>     @	@   <�D�?��ƀ�7>     �	@   h)P�?R`D�OG>     �	@   �T[�?9%� ��K>      
@   �Mf�?��/�<>     @
@   �q�?�Ò��?>     �
@   �{�?4��2G<>     �
@   L��?Â���|/>      @   �Y��?���s�
@>     @@   �k��?��Ò�a@>     �@   XS��?x(3��u8>     �@   ���?v�O,ib>      @   ȥ��?�&L͒C>     @@   ���?��}��L>     �@   �X��?Lo����>     �@   �x��?-�Ϡ�9>      @   �s��?6FID?9>     @@   8J��?����gsL>     �@   d���?��y>     �@   ���?>�&�09C>      @   ����?
��<�A>     @@   (J�?I�V	C>     �@   `w�?��^@�N>     �@   ���?�#��%�@>      @   �s�? �M�K>     @@    D'�?ή�Q��->     �@   ��.�?9!���G>     �@   ��6�?.����1>      @   >�?.1�NcB>      @   �cE�?�sǔ�1>     @@   L�L�?�n�HN>     `@   H�S�?�W��$>     �@   8�Z�?
Ȃ�q�;>     �@   ��a�?N�/�[7>     �@   (�h�?�=�mC>     �@   0oo�?�H75M>      @   Hv�?P��.�#>      @   �|�?�G���7>     @@   �*��?�#4��2I>     `@   ����?o���oJ>     �@   ����?���-��#>     �@   ���?�h��%F>     �@   @��?R�x^D>     �@   PP��?�� s�@>      @   4L��?P�_!
�#>      @   4��?��:#�G>     @@   L��?qg�:&J>     `@   Hɹ�?5L$.��4>     �@   \w��?!�1�C>     �@   ���?���[<>     �@   D���?��<���=     �@   ���?��
~���=      @   �y��?������B>      @   ����?�~.���4>     @@   h��?��u�|�8>     `@   �E��?A8yL;>     �@   �h��?��41��C>     �@   �{��?-���+oF>     �@   $��?x���O>     �@   s��?�՝m�T2>      @   �W��?����=>      @   �-�?î�\�=>     @@   ��?���\=�=     `@   ��?j\&">     �@   �X�?��1�D>>     �@   ���?�#O#`�I>     �@   ��?�}���0>     �@   ��?���F\IE>      @   t{#�?��ׯ,B>      @   0�'�?�E� ]�$>     @@   ,>,�?��ކ?5>     `@   ��0�?��iIqE>     �@   ��4�?�ha�;>     �@   �9�?��A���D>     �@   �.=�?̤KF�w�=     �@   DMA�?�����=      @   `E�?ap�I0�H>      @   �gI�?��:���->     @@   �cM�?��%Q>     `@   @UQ�?Ly5ښoE>     �@   �;U�?v�g�0�/>     �@   �Y�?jv�U�G>     �@   �\�?�����yK>     �@   ,�`�?A%My��>      @   md�?���H>      @    h�?�p���M>     @@   0�k�?k��}<>     `@   �ho�?����f7O>     �@   ��r�?���}�O>     �@    �v�?+��i�I>     �@   @z�?�b�B'=>>     �@   `�}�?Z����M>      @   ����?1�����M>      @   �a��?R�~���=     @@   t���?QNT	��B>     `@   x��?�W3c�L>     �@   g��?�+(����=     �@   D���?q���J�K>     �@   L��?� ;,*>     �@   8!��?������D>      @   ,O��?� ����E>      @   Du��?��in]D>     @@   ����?%����3F>     `@   P���?^��F"VM>     �@   ����?�}�30}->     �@   @���?�~F	y�;>     �@   ����?l	R(>     �@   躰�?��\�7`>      @    ���?�dg���;>      @   ���?�;Sv�@E>     @@   <|��?�����M>     `@   �Y��?|}�;�2>     �@   ,0��?�<v��G>     �@   $ ��?̯�/p�">     �@   ����?���\(0>     �@   |���?[s$���F>      @   I��?�d�ӔV>      @   T���?���0)LK>     @@   h���?�)�5G�5>     `@   XY��?�|��zJ>     �@   @���?W�޾�L?>     �@   0���?����6:>     �@   <3��?��Q���B>     �@   x���?7o��/�M>      @   �Q��?�Kc�Z�0>      @   ����?�z-�A5>     @@   Z��?"B�DcI>     `@   ����?��`I�.>     �@    L��?L�d�%>     �@   ���?"�l"w �=     �@   �(��?�?��!>     �@   ���?��j^�J>      @   8���? ϞH��0>      @   LL��?���%�C>     @@   T���?��J�+N>     `@   d���?;l�>�0>     �@   �B��?�^{v�@>     �@   Ȋ��?�@Y˕B>     �@   @� �?T�l���0>     �@   ��?w4n4>      @    G�?�oN�=�;>      @   h|�?�L�{�/>     @@   <�	�?B�nu5>     `@   ���?���`�,+>     �@   d�?����5>     �@   �$�?l��  >     �@   �C�?~+^��M>     �@   �^�?�PK�QD >      @   ,u�?^{�#tF>      @   |��?�^4K�� >     @@   ���?��4�O
>>     `@   ���?XEړ� J>     �@   ���?(�gԹ�,>     �@   �� �?43-spF>     �@   ��"�?P`E5�+*>     �@   ��$�?=�QQ�D>       @-DT�!�?\3&��<( n u l l )     (null)         EEE50 P    ( 8PX 700WP        `h````  xpxxxx                                                                                                                                                                                                                                                                                                ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ 1#QNAN  1#INF   1#IND   1#SNAN  C O N O U T $   ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp           H                                                           �1 "   RSDS^�.lkeE��6s*�.�   C:\Program Files\MAXON\CINEMA 4D R12\plugins\Maze Trace\obj\cinema4dsdk_Win32_Release.pdb              ,4     0        ����    @                0d           t�4     0       ����    @   d           ���    80       ����    @   �P0        ����    @   �            �               (��    h0       ����    @               �0X           h|(��    �0       ����    @   X            �0�           ��(��    �0       ����    @   �            P0�            �0            $ ,     �0        ����    @                �0\            l x 4    �0       ����    @   \             �0�            � �     �0        ����    @   �             1�             !!    1        ����    @   �             418!           H!T!4    41       ����    @   8!            X1�!           �!�!    X1        ����    @   �!            �1�!           �!�!    �1        ����    @   �!�� @ �h                     ����    ����    ����    ��    ����    ����    ������	�    ����    ����    ����    ;    ����    ����    ����    #�    ����    ����    ����    ������    �����    ����    ����    ������    ������    ����    ����    �    ����    ����    ����    X	    ����    ����    ����    *    ����    ����    ����    �    ����    ����    ����    g    ����    ����    ����    �    ����    ����    �����$�$    ����    ����    ����;&N&    ����    ����    ����040    ����    ����    ����    �k    ����    ����    ����    �s    ����    ����    ����    |    ����    ����    ����    E~    ����    ����    ����    �        �����    ����    ����    0�    ����    ����    ����    	�    ����    ����    ����    փ<%         �*  �                     @& P& `& v& �& �& �& �& �& �& �& �& 
' ' &' 0' H' \' l' �' �' �' �' �' �' �' ( ( 4( N( d( ~( �( �( �( �( �( �(  ) ) () D) b) v) �) �) �) �) �) �) �) �) * * &* <* N* `* p* �* �* �* �* �*     � DecodePointer � EncodePointer �GetCurrentThreadId  �GetCommandLineA �HeapAlloc GetLastError  �HeapFree  %WriteFile dGetStdHandle  GetModuleFileNameW  IsProcessorFeaturePresent �TlsAlloc  �TlsGetValue �TlsSetValue �TlsFree �InterlockedIncrement  GetModuleHandleW  sSetLastError  �InterlockedDecrement  EGetProcAddress  �Sleep ExitProcess oSetHandleCount  �InitializeCriticalSectionAndSpinCount �GetFileType cGetStartupInfoW � DeleteCriticalSection GetModuleFileNameA  aFreeEnvironmentStringsW WideCharToMultiByte �GetEnvironmentStringsW  �HeapCreate  �HeapDestroy �QueryPerformanceCounter �GetTickCount  �GetCurrentProcessId yGetSystemTimeAsFileTime �HeapSize  �TerminateProcess  �GetCurrentProcess �UnhandledExceptionFilter  �SetUnhandledExceptionFilter  IsDebuggerPresent rGetCPInfo hGetACP  7GetOEMCP  
IsValidCodePage 9LeaveCriticalSection  � EnterCriticalSection  RtlUnwind ?LoadLibraryW  �HeapReAlloc �RaiseException  -LCMapStringW  gMultiByteToWideChar iGetStringTypeW  fSetFilePointer  �GetConsoleCP  �GetConsoleMode  �SetStdHandle  $WriteConsoleW � CreateFileW R CloseHandle WFlushFileBuffers  KERNEL32.dll      Gl�Q    +          + + +  � "+   cinema4dsdk.cdl c4d_main                                                                                                                                                                                                                      ��    .?AVGeSortAndSearch@@   ��    .?AVSorter@@    ��    .?AVNodeData@@  ��    .?AVBaseData@@  ��    .?AVObjectData@@    ��    .?AVPointGeneratorData@@    ��    .?AVTSPData@@   ��    .?AVNeighbor@@  ��    .?AVDisjointNgonMesh@@  ��    .?AVGeToolNode2D@@  ��    .?AVGeToolDynArray@@    ��    .?AVGeToolDynArraySort@@    ��    .?AVGeToolList2D@@  u�  s�      sqrt    ��    .?AVtype_info@@ asin            acos            cos             sin             atan            log N�@���D    OOOOOOOOOO           ��������    �����
                                                                                           	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                 ?                                                                                                                                                                                                                                                                                                                                                  abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                      4�  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��    ����C   ����������������x�p�d�X�P�D�@�<�8�4�0�,�(�$� ����� �����0�����������������������x�	         p�h�`�X�P�H�@�0� ��������������������������|�t�l�d�T�@�4�(����� ���������������h�T�                                                                                           $9            $9            $9            $9            $9                              �=        H�P(9�:                                                                                                                                                                                                                                                                                      �&         ��   ��   ��   ��   ��   ��!   ��   ��   |�   l�   ��   ��   P�   L�    H�   d�   \�   ��   T�   ��   ��   x�   p�   h�"   d�#   `�$   \�%   T�&   H�      �      ���������              �       �D        � 0     ��    .   .   �=QQQQQQQQQ�=QQQQQQQ�=HJL   ���5      @   �  �   ����                      �            @Q    @Q                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                .                   �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
    ����                                               |   �0�0T1g12+2=2V2�4�45"535E5N5b5{5�5�5�5�566~6�6�6�68�9:$:D:L<t<�<�<�<�<�<�<=(=T=f=�=�=
>K>d>�>�>?o?�?�?�?�?�?    X   00#01D1]1�1e2�23�3�34$4m4�4	56)6=6 77�7�7[9d9�9�:�:�;�;�;==9=�>�>�?�?�? 0  �   �0�0�0�1�1�3�344(4T4j4|4�4�4�4�4�4585K5�5�56w6�6�647F7[7a7�7�7�7�7!838D8V8�9�9�9�9�9:=;n;�;�;�;<D<�<�<=�=�=~>�>�>�?�? @  |   H0M0�1�12�3�334=4Y4�5�5�5�6�6�6�7�7�7�7$8D8a8�8�8I9e9�9�9I:e:�:�:;,;H;d;�;�;<%<�<�<<=a=�=�=>$>D>d>q>�>�>�>?$?   P  d   �8�8�8.9d9x9�9�9�9":::v:�:�:�: ;1;�; <<I<S<d<�<�<�<�<=K=\=�=�=�=�=>>>>>F>W>k>>�>�>
?�? `  �   h3l3p3t3x3|394P4a4n5�5�6�6�6�6�6%7+7O7t7�7�7�7�7�788?8d8�8�8�8�9�9	::":y:�:;L;P;T;X;\;<<A<T<�<�<�<�<=�=�=�=4>d>�>�>?$?D?a?�?�?�? p  8  0$0Y01$1D1{1�1�12�2�2�23>3Y3�3�3�3'4[4�4�4�4�4�4
5$515>5V5i5{5�5�5�5�5�5�56(6D6U6h6�6�6�6�6�6�6�67767T7f7�7�7�7�7�7�7�7 868R8c8v8�8�8�8�8�8�899(9F9d9v9�9�9�9�9�9�9:0:F:b:t:�:�:�:�:�: ;;$;D;R;_;w;�;�;�;�;�;�;<<2<H<d<v<�<�<�<�<�<==&=/=M=n=�=�=�=�=�=�=>">>>O>b>�>�>�>2?:?D?V?`?{?�?�?�?�?�?   �  �   /0Q0f0�0�0�0�0�01e1w1�1�1�1�1242T2h2z2�2�2�233�3�3�3A4�4�4�4�4�45$5D5a5t5�5�5�5*7<7N7�7P8W8^8e8l8s8z8�8�8�8�8�8�8�8�8�8�8:-:Z:y:�:�:�:�;�;�;�<>>>!>+>5>?>T>�>�>�>�>�>�?�?�? �  �   00D0t0�0�0�0141T1�1�1�1242T2t2�2�2�2�23&3A3T3q3�3�3�3�3�34Q4a4t4�4�4�4545Q5a5q5�5�5�5�56$6D6o6�6�6�6�67$7D7d7�7�7�7�748Z8�8�8�8�89$9D9d9�9�9�9�9':g:�:�:#;d;�;�;�;$<Q<q<�<�<�<�<==4=T=t=�=�=�=�=6>T>q>�>�>�>�>$?D?d?�?�?�?�? �    020F0V0�0�0�0�01$1P1d1t1�1�1�12*2]2k2~2�2�2�2�2�23.3B3R3t3�3�3�3�34(4T4l4�4�4�4�4 55'565d5|5�5�5�5�56)676F6t6�6�6�6�677T7}7�7�7�7�7�748T8t8�8�8�89$9D9d9�9�9�9�9�9$:D:d:�:�:�:�:;$;D;d;�;�;�;�;�;<!<1<T<i<{<�<�<�<�<�<�<�<$=T=t=�=�=�=>4>Q>t>�>�>�>?D?t?�?�?   �  �   0R0q0�0�0�0�0$1Q1q1�1�1�1�1$2T2�2�2�2�2343T3�3�3�3�3�3!404T4�45A5T5t5�5�5�5!6A6q6�6�6�67!7D7�7�7�7848d8�8�8�8:9{9�9�9�9:4:d:�:�:�:�:�:;J;d;�;�;<*<t<�<�<p=�=>%>:>]>�>�>�>?6?_?�?�?�?   �  �   0H0y0 1D1T1�1�1�1	232G2e2�2�2�2�23D3d3�3�3�3�34a4�4�4�45!5D5d5�5�5�5$6q6�6�6�6�6?7^7z7�7�7�7(8C8q8�8�8�8�89&9V9x9�9�9�9�9:3:H:�:�:�:�:;+;K;`;|;;<N<�<�<�<�<=d=w? �  �   282�2�2�2�23T3o3$5(5,505k5p5�5�5�566D6d6�6�6�6�6$767d7�7�7�7�788A8d8�8�8�8�89$9Q9d9�9�9�9:1:Q:t:�:�:�:!;A;d;�;�;�;<4<T<t<�<�<�<�<=4=T=q=�=�=�=�=>n>�>�>?G?�?�?   �  �   !0�0�0�0X1z1�12.2F2�2�2�2s3�3�3�34d45,5T5�5�5$6�6�6�6n7�7�78�8�8979�9�9:7:�:�:s;�;�;><^<s<�<=#=w=�=<>�>�>�>?!?4?d?�?�?�?�?   �    040q0�0�0�0�0141g1�1�1�12>2W2k2�2�2�2313T3q3�3�3N4S4X4]44�4�4�45$5D5d5�5�5�5646Q6a6q6�6�67@7n7�7�78>8q8�8�8�8�8�89%939T9e9s9�9�9�9�9:!:1:T:l:�:�:�:�:�: ;;;0;T;l;�;�;�;�;�;�;
<<+<=<a<q<�<�<�<�<=4=F=T=g=�=�=�=>$>A>T>t>�>�>�>??4?T?t?�?�?�?�?�?     (  0$0D0d0�0�0�0�01'1X1j11�1�1�12D2o2�2�2�23$3D3d3�3�3�3�34!444d4�4�4�4�4�455-5;5J5\5�5�5�5�5�56$6Q6a6q6�6�6�6�6�6�6�677,7T7t7�7�7�7�7848T8t8�8�8�8�89)9E9]9w9�9�9�9�9:4:T:t:�:�:�:�:�:�:;";1;A;S;t;�;�;�;�;�;<"<7<Q<b<�<�<�<�<�<�<1=D=t=�=�=�=�=�=>$>D>d>�>�>�>�>?$?D?d?�?�?�?�?  �   0$0D0d0�0�0�0 1$1D1d1�1�1�1�12$2D2d2�2�2�2�23$3D3d3�3�3�3�34$4D4a4t4�4�4�4�45!515A5T5t5�5�5�5�56$6D6^6f6}6�6�67!747G7h7�7d8�8�8�859r9�9�9E:u:�:�:;a;�;�;%<e<�<�<=U=�=�=>e>�>�>?E?�?�?�?     �   50�0�01E1�1�1�1�1�12e2�2�2"3e3�3�3B4�4�4�4	55@5E5m5�5�5�5	6E6i6�6�6%7I7r7�7�78/8h8�8�8�8989v9�9�9$:A:d:�:�:�:;A;T;�;�;�;�;<4<S<f<�<�<�<=1=D=t=�=�=�=>T>�>�>�>�>$?D?a?�?�?�?�?   0 �   040f0{0�0!141d1�1�1�1�3�3�3�3�5�5�5$6T6t6�6�6�6�67D7t7�7�7�7�78!8D8a8t8�8�8�9�9J:O:�:�;�;�;�<�<�<=Q=[=�=�=>4>�>�>$?d?�?�?�?�?   @ �   0$0D0d0�0�0�0�0$1D1q1�1�1�12A2d2�2�2�2!3A3a3�3�3�3�34!4A4a4�4�4�4�45!5A5a5�5�5�5�56$6D6a6�6�6�6�6747T7q7�7�7�78�8�8   P T   �4�4�4%5e5�5�556u6�6�67U7�7�78E8�8�8�8"9R9�9�9�95:�:�:;U;�;�;%<�<�<�>�>�? ` �   �1X2\2`2d2h2K3Y3x3�34&4K4S45 5Q5_5�5�5�6�6�67p7~7�7�7�8�8�89$9D9d9�9�9�9�9�9::$:A:T:t:�:�:�:�:;4;Q;t;�;�;�;<$<D<d<�<�<�<==$=D=d=�=�=�=�=>>D>o>�>�>�>??,?Q?d?�?�?�?�?�?�?   p |   �0�021e1�152u2�23E3�3�3"4R4�4�4%5e5�5�5B6u6�6"7R7�7�7�7"8U8�8�8(9<9L9j9�9�9:e:�:�:E;�;�;5<�<�<=R=�=�=">h>�>"?h?�? � t   "0e0�01U1�1�1B2�23�34E4�4�45U5�5�556�6�6%7r7�78U8�89U9�9�9�9:U:�:�:%;u;�;<e<�<=v=�=>E>�>�>?U?�?�? � |   N0u0�0 1M1t1�12o2�2�2L3�3 4444A4G4s4z4�4�4�4�45$5(5,5054585A5d5�5646�6�6X7i7�:=;M;�<�<E=t={=�=�=�=�==>�>�>?�?�? � �   �061�1�1�1�12*3�3<4d4D5d5�5�5�5!6D6t6�6�6�6$7T7�7�7=8D8K8R8Y8`8g8n8x8�8�8�8�8�8�8�8�8�8�8�8�8�8959m9~9�9D:�:�;�;�;�;�;�;�;�;�;�;�;�;<<<<<< <�<�<�<�<�<�<2=N= >�>�>�>�>�>�>�>�>???]?d?h?l?p?t?x?|?�?�?�?�?�?�?   �   B0M0h0o0t0x0|0�0�0�0 11111111f1l1p1t1x1�1�122?2W2_2h2�2�2�2�2�2(3D3\3�3�3P44�4�4�4�4�45R5�5�56.696K6b6�6%777~7�7�7�7�7Y8g8y8�8�8�8�8�8"9�9�9�9�9�9�9�9:Z:s:�:;;";B;�;�;�;<'<=<O<b<�<='=4=d=�=�=�=�=�=�=9>>>G>V>y>~>�>�>�>*?\?t?{?�?�?�?�?�?�?�? � p   0000000 0j0p0t0x0|0�0�011111=1g1�1�1�1�1�1�1�1�1�122222�2�2�2�2i5�56e;&<�=�=�=)>�>8?�? � H  k0l1|1�1�1�1�1�1�1�1�2�233d3|3�3�3�3�3�3�3�34D4a4�4�4555�6�6�6�6�67777(7.767<7H7N7[7e7k7u7�7�7�788B8H8N8d8|8�89?9I9�9�9�9�9�9�9�9:::(:6:@:F:\:a:i:o:v:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:	;;;;$;);1;6;=;L;Q;W;`;�;�;�;�;�;�;<&<2<k<t<�<�<�<�<�<�<I=Q=d=o=t=�=�=�=�=�=�=�=�=>	>>>0>i>s>�>�>�>�>�>k?�?�?�? � �   00"0i0s0�0�0�0�0(1:1h1�1�1�1�1�1�12=2G2�2�2�2�2�2y4�4�4�4�4�45515Y5�5�5�5�5�5�566(6.646A6^6�6�7�7�7�78�9�9�9�9�9�9�9#:+:A:]:�:�:�:�:�:�:�:2;:;F;�;�;�;�;<u<�<�<�<�<===�=�=�=>>'>c>�>�>�>�> �   000�0�0�0$111]1e1�1�1T2l2�2�2�2�2)353=3I3�3�3�3�3�3484�5�5�5�5)656E6Q6n6t6�6�6�6�6~7�7�7�788$898^8�8�8*9@9P9z9�9�9�9�98:q:z:�:�:�:�:�:�:�:;=;X;_;h;q;z;�;�;�;�;�;�; <<<<<<<< <$<(<,<0<E<�<:=B=V=`=~=�=�=�=�=�=�=>>>(>4>@>t>~>�>�>�>�>�>�>?? ?,?d?s?{?�?�?�?�?�?�?   �   90A0I0Q0o0w0�0�0�011h1�1�1�1�1�1�1�23Q3�3�3�3�34�4�4o5u5{5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 6	66 6%656:6@6F6\6c6�6<7S7�8�899%939<9F9z9�9�9�9�9�9�9 :U:h:�:�:>;�;�;A<M<`<r<�<�<�<�<�<�<�<�<===<=e=v=�=�=%>m>�>�?�?  �   *0D0U0�0�0�0�1�1�1
222$2�2�2�34�4�7�9�:�:;; ;7;E;K;n;u;�;�;�;�;�;�;(<|<�<�<�<�=>>>>*>Y>_>g>�>�>�>�>�>�>?
??y?�?�?   �   030>0D0T0Y0j0r0x0�0�0�0�0�0�0�0�0�0�0�01.1H1J3Q3W3�3�3�3O4U4a4�4�4�4�4555�5�5�5�566 9f:�:�:�:�:";+<�<�<1=�=�?�?�?�?�? 0 L   	090�0�0M1X1�1�1�2�2�3�4�4�4>5M5h5}8s9;J;v;�;{=�?�?�?�?�?�?�?�?�?   @ X   0M0�0�102S2�2�6�6�677E7W7i7{7�7�7�7�7�7�7�78899�9�:�:i;J<�<�<�=�=�=9>P>�>? P L   0	0�0�13292�2�2�2�3�3�3^4727~:�:�:�:�:�:�:�:�:�:�:�:�:y;�;�;�;<C< ` 0   J6�899�9�9�9�:�:;!;];�;<w<=:=*>S>�> p �   0�0�1�12L2k23:3b3�3D4g4y44�4�4�4�4�4�4�4�4 5$565D5Y5c5�5�5�5�5�5'6T6_6s7�7�:�:�:�:<;d;};�;�;�;�;,<:<H<U<t<=�=�=�=�=>>>&>?$?/?R?�?   � <   3090>0D0U0�0>1h1�1�1�1�2�2�2�2 3R3z34!424:4D4V4`4{4 � �   1111 1$10141�1�1(2,2024282<2@2D2H2L2P2T2X2\2`2d2h2l2p2t2x2|2�2�2�2�2�2�2�2�2�2�2�2`3d3h3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3d5h5�5�5�5�5�54787�7�7�7�7�7�7�7�7�7 � 4   111$1,141<1D1L1T1\1d1l1t1|1�1�1�1�1�1�1�1 � �   :0>0B0F0L0P0H9L9P9T9X9\9`9d9h9l9p9t9x9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 :::::::: :$:(:,:0:4:8:<:@:D:H:L:P:T:X:\:`:d:h:l:p:t:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:    h   �=�=(>,>4>L>\>`>p>t>x>�>�>�>�>�>�>�>�>�>�> ???? ?(?@?P?T?d?h?l?p?t?|?�?�?�?�?�?�?�?�?�?�?�?�?   �   00 0$0,0D0T0X0h0l0p0x0�0�0�0�0�0�0�0�0�0�0 11 10141D1H1L1T1l1|1�1�1�1�1�1�1�1�1�1�1�182T2X2x2�2�2�2�2�23(3H3h3�3�3�3�3�3�344(4H4h4�4�4�4�4�45 0 l   0 080P0h0�0�0�0�0�0141X1�1 22222222 2$2(8(9,9094989<9@9D9H9L9P9T9X9\9`9d9h9l9p9t9x9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 :::::::: :$:(:,:0:4:8:<:@:D:H:L:P:T:X:\:`:d:h:l:p:t:x:|:�:�:�:�:�:;;(;L;X;\;`;d;h;�<�<�<�<�<�<�<�<�<�<�<�<�<====$=,=4=<=D=L=T=\=d=l=t=|=�=�=�=�=�=�=�=�=�=�=�=�=>>>>>> >$>(>,>0>4>�>�>                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  